magic
tech sky130A
magscale 1 2
timestamp 1641609411
<< nwell >>
rect -636 0 1036 626
<< pwell >>
rect -626 -644 1026 -432
<< psubdiff >>
rect -600 -521 1000 -458
rect -600 -555 -531 -521
rect -497 -555 -463 -521
rect -429 -555 -395 -521
rect -361 -555 -327 -521
rect -293 -555 -259 -521
rect -225 -555 -191 -521
rect -157 -555 -123 -521
rect -89 -555 -55 -521
rect -21 -555 13 -521
rect 47 -555 81 -521
rect 115 -555 149 -521
rect 183 -555 217 -521
rect 251 -555 285 -521
rect 319 -555 353 -521
rect 387 -555 421 -521
rect 455 -555 489 -521
rect 523 -555 557 -521
rect 591 -555 625 -521
rect 659 -555 693 -521
rect 727 -555 761 -521
rect 795 -555 829 -521
rect 863 -555 897 -521
rect 931 -555 1000 -521
rect -600 -618 1000 -555
<< nsubdiff >>
rect -600 525 1000 588
rect -600 491 -531 525
rect -497 491 -463 525
rect -429 491 -395 525
rect -361 491 -327 525
rect -293 491 -259 525
rect -225 491 -191 525
rect -157 491 -123 525
rect -89 491 -55 525
rect -21 491 13 525
rect 47 491 81 525
rect 115 491 149 525
rect 183 491 217 525
rect 251 491 285 525
rect 319 491 353 525
rect 387 491 421 525
rect 455 491 489 525
rect 523 491 557 525
rect 591 491 625 525
rect 659 491 693 525
rect 727 491 761 525
rect 795 491 829 525
rect 863 491 897 525
rect 931 491 1000 525
rect -600 428 1000 491
<< psubdiffcont >>
rect -531 -555 -497 -521
rect -463 -555 -429 -521
rect -395 -555 -361 -521
rect -327 -555 -293 -521
rect -259 -555 -225 -521
rect -191 -555 -157 -521
rect -123 -555 -89 -521
rect -55 -555 -21 -521
rect 13 -555 47 -521
rect 81 -555 115 -521
rect 149 -555 183 -521
rect 217 -555 251 -521
rect 285 -555 319 -521
rect 353 -555 387 -521
rect 421 -555 455 -521
rect 489 -555 523 -521
rect 557 -555 591 -521
rect 625 -555 659 -521
rect 693 -555 727 -521
rect 761 -555 795 -521
rect 829 -555 863 -521
rect 897 -555 931 -521
<< nsubdiffcont >>
rect -531 491 -497 525
rect -463 491 -429 525
rect -395 491 -361 525
rect -327 491 -293 525
rect -259 491 -225 525
rect -191 491 -157 525
rect -123 491 -89 525
rect -55 491 -21 525
rect 13 491 47 525
rect 81 491 115 525
rect 149 491 183 525
rect 217 491 251 525
rect 285 491 319 525
rect 353 491 387 525
rect 421 491 455 525
rect 489 491 523 525
rect 557 491 591 525
rect 625 491 659 525
rect 693 491 727 525
rect 761 491 795 525
rect 829 491 863 525
rect 897 491 931 525
<< poly >>
rect -506 -42 -476 36
rect 94 -42 124 36
rect 294 -42 324 36
rect 894 -42 924 36
<< locali >>
rect -576 525 976 566
rect -576 491 -537 525
rect -497 491 -465 525
rect -429 491 -395 525
rect -359 491 -327 525
rect -287 491 -259 525
rect -215 491 -191 525
rect -143 491 -123 525
rect -71 491 -55 525
rect 1 491 13 525
rect 73 491 81 525
rect 145 491 149 525
rect 251 491 255 525
rect 319 491 327 525
rect 387 491 399 525
rect 455 491 471 525
rect 523 491 543 525
rect 591 491 615 525
rect 659 491 687 525
rect 727 491 759 525
rect 795 491 829 525
rect 865 491 897 525
rect 937 491 976 525
rect -576 452 976 491
rect 94 382 420 416
rect -632 310 -458 344
rect 94 342 128 382
rect -632 14 -598 310
rect 386 266 420 382
rect 370 232 420 266
rect 648 14 682 58
rect -632 -20 682 14
rect -576 -521 976 -482
rect -576 -555 -537 -521
rect -497 -555 -465 -521
rect -429 -555 -395 -521
rect -359 -555 -327 -521
rect -287 -555 -259 -521
rect -215 -555 -191 -521
rect -143 -555 -123 -521
rect -71 -555 -55 -521
rect 1 -555 13 -521
rect 73 -555 81 -521
rect 145 -555 149 -521
rect 251 -555 255 -521
rect 319 -555 327 -521
rect 387 -555 399 -521
rect 455 -555 471 -521
rect 523 -555 543 -521
rect 591 -555 615 -521
rect 659 -555 687 -521
rect 727 -555 759 -521
rect 795 -555 829 -521
rect 865 -555 897 -521
rect 937 -555 976 -521
rect -576 -594 976 -555
<< viali >>
rect -537 491 -531 525
rect -531 491 -503 525
rect -465 491 -463 525
rect -463 491 -431 525
rect -393 491 -361 525
rect -361 491 -359 525
rect -321 491 -293 525
rect -293 491 -287 525
rect -249 491 -225 525
rect -225 491 -215 525
rect -177 491 -157 525
rect -157 491 -143 525
rect -105 491 -89 525
rect -89 491 -71 525
rect -33 491 -21 525
rect -21 491 1 525
rect 39 491 47 525
rect 47 491 73 525
rect 111 491 115 525
rect 115 491 145 525
rect 183 491 217 525
rect 255 491 285 525
rect 285 491 289 525
rect 327 491 353 525
rect 353 491 361 525
rect 399 491 421 525
rect 421 491 433 525
rect 471 491 489 525
rect 489 491 505 525
rect 543 491 557 525
rect 557 491 577 525
rect 615 491 625 525
rect 625 491 649 525
rect 687 491 693 525
rect 693 491 721 525
rect 759 491 761 525
rect 761 491 793 525
rect 831 491 863 525
rect 863 491 865 525
rect 903 491 931 525
rect 931 491 937 525
rect -537 -555 -531 -521
rect -531 -555 -503 -521
rect -465 -555 -463 -521
rect -463 -555 -431 -521
rect -393 -555 -361 -521
rect -361 -555 -359 -521
rect -321 -555 -293 -521
rect -293 -555 -287 -521
rect -249 -555 -225 -521
rect -225 -555 -215 -521
rect -177 -555 -157 -521
rect -157 -555 -143 -521
rect -105 -555 -89 -521
rect -89 -555 -71 -521
rect -33 -555 -21 -521
rect -21 -555 1 -521
rect 39 -555 47 -521
rect 47 -555 73 -521
rect 111 -555 115 -521
rect 115 -555 145 -521
rect 183 -555 217 -521
rect 255 -555 285 -521
rect 285 -555 289 -521
rect 327 -555 353 -521
rect 353 -555 361 -521
rect 399 -555 421 -521
rect 421 -555 433 -521
rect 471 -555 489 -521
rect 489 -555 505 -521
rect 543 -555 557 -521
rect 557 -555 577 -521
rect 615 -555 625 -521
rect 625 -555 649 -521
rect 687 -555 693 -521
rect 693 -555 721 -521
rect 759 -555 761 -521
rect 761 -555 793 -521
rect 831 -555 863 -521
rect 863 -555 865 -521
rect 903 -555 931 -521
rect 931 -555 937 -521
<< metal1 >>
rect -592 536 1010 566
rect -592 525 183 536
rect 235 525 1010 536
rect -592 491 -537 525
rect -503 491 -465 525
rect -431 491 -393 525
rect -359 491 -321 525
rect -287 491 -249 525
rect -215 491 -177 525
rect -143 491 -105 525
rect -71 491 -33 525
rect 1 491 39 525
rect 73 491 111 525
rect 145 491 183 525
rect 235 491 255 525
rect 289 491 327 525
rect 361 491 399 525
rect 433 491 471 525
rect 505 491 543 525
rect 577 491 615 525
rect 649 491 687 525
rect 721 491 759 525
rect 793 491 831 525
rect 865 491 903 525
rect 937 491 1010 525
rect -592 484 183 491
rect 235 484 1010 491
rect -592 452 1010 484
rect -592 62 -558 452
rect -8 378 326 412
rect -524 292 -458 360
rect -326 352 -256 362
rect -326 300 -317 352
rect -265 300 -256 352
rect -326 290 -256 300
rect -8 262 26 378
rect 292 350 326 378
rect 674 352 744 362
rect 76 294 142 350
rect 276 294 342 350
rect 674 300 683 352
rect 735 300 744 352
rect 674 290 744 300
rect 876 292 942 360
rect -424 62 -358 262
rect -8 228 42 262
rect 176 232 242 262
rect 176 180 183 232
rect 235 180 242 232
rect 176 62 242 180
rect 776 62 842 262
rect 976 62 1010 452
rect -564 20 -498 26
rect -270 20 -224 62
rect -564 19 -224 20
rect -564 -33 -557 19
rect -505 -26 -224 19
rect -505 -33 -498 -26
rect -564 -40 -498 -33
rect -558 -68 -512 -40
rect 42 -68 88 62
rect 330 -68 376 62
rect 642 20 688 62
rect 916 20 982 26
rect 642 19 982 20
rect 642 -26 923 19
rect 916 -33 923 -26
rect 975 -33 982 19
rect 916 -40 982 -33
rect 930 -68 976 -40
rect -430 -268 -358 -68
rect -224 -268 -158 -68
rect -24 -268 42 -68
rect -416 -482 -358 -268
rect -324 -306 -258 -300
rect -324 -358 -316 -306
rect -264 -358 -258 -306
rect -324 -364 -258 -358
rect -124 -307 -58 -300
rect -124 -359 -117 -307
rect -65 -359 -58 -307
rect -124 -366 -58 -359
rect 130 -482 288 -68
rect 376 -268 442 -68
rect 576 -268 642 -68
rect 776 -268 842 -68
rect 476 -307 544 -300
rect 476 -356 485 -307
rect 478 -359 485 -356
rect 537 -359 544 -307
rect 478 -366 544 -359
rect 676 -306 742 -300
rect 676 -358 684 -306
rect 736 -358 742 -306
rect 676 -364 742 -358
rect 776 -482 834 -268
rect -576 -521 976 -482
rect -576 -555 -537 -521
rect -503 -555 -465 -521
rect -431 -555 -393 -521
rect -359 -555 -321 -521
rect -287 -555 -249 -521
rect -215 -555 -177 -521
rect -143 -555 -105 -521
rect -71 -555 -33 -521
rect 1 -555 39 -521
rect 73 -555 111 -521
rect 145 -555 183 -521
rect 217 -555 255 -521
rect 289 -555 327 -521
rect 361 -555 399 -521
rect 433 -555 471 -521
rect 505 -555 543 -521
rect 577 -555 615 -521
rect 649 -555 687 -521
rect 721 -555 759 -521
rect 793 -555 831 -521
rect 865 -555 903 -521
rect 937 -555 976 -521
rect -576 -594 976 -555
<< via1 >>
rect 183 525 235 536
rect 183 491 217 525
rect 217 491 235 525
rect 183 484 235 491
rect -317 300 -265 352
rect 683 300 735 352
rect 183 180 235 232
rect -557 -33 -505 19
rect 923 -33 975 19
rect -316 -358 -264 -306
rect -117 -359 -65 -307
rect 485 -359 537 -307
rect 684 -358 736 -306
<< metal2 >>
rect 176 536 242 542
rect 176 484 183 536
rect 235 484 242 536
rect -326 352 -256 362
rect -326 300 -317 352
rect -265 300 -256 352
rect -326 110 -256 300
rect 176 232 242 484
rect 176 180 183 232
rect 235 180 242 232
rect 176 174 242 180
rect 674 352 744 362
rect 674 300 683 352
rect 735 300 744 352
rect 674 110 744 300
rect -326 40 744 110
rect -564 19 -498 26
rect -564 -33 -557 19
rect -505 -33 -498 19
rect -564 -40 -498 -33
rect -564 -106 -58 -40
rect -322 -306 -258 -300
rect -322 -358 -316 -306
rect -264 -358 -258 -306
rect -322 -420 -258 -358
rect -124 -307 -58 -106
rect -124 -359 -117 -307
rect -65 -359 -58 -307
rect -124 -366 -58 -359
rect 174 -420 244 40
rect 916 19 982 26
rect 916 -33 923 19
rect 975 -33 982 19
rect 916 -40 982 -33
rect 478 -106 982 -40
rect 478 -307 544 -106
rect 478 -359 485 -307
rect 537 -359 544 -307
rect 478 -366 544 -359
rect 678 -306 742 -300
rect 678 -358 684 -306
rect 736 -358 742 -306
rect 678 -380 742 -358
rect 676 -420 742 -380
rect -322 -484 742 -420
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_0
timestamp 1641609411
transform 1 0 909 0 1 -168
box -99 -126 99 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_1
timestamp 1641609411
transform 1 0 309 0 1 -168
box -99 -126 99 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_2
timestamp 1641609411
transform 1 0 109 0 1 -168
box -99 -126 99 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_3
timestamp 1641609411
transform 1 0 -491 0 1 -168
box -99 -126 99 126
use sky130_fd_pr__nfet_01v8_59MFY5  sky130_fd_pr__nfet_01v8_59MFY5_0
timestamp 1641609411
transform 1 0 709 0 1 -199
box -99 -157 99 157
use sky130_fd_pr__nfet_01v8_59MFY5  sky130_fd_pr__nfet_01v8_59MFY5_1
timestamp 1641609411
transform 1 0 509 0 1 -199
box -99 -157 99 157
use sky130_fd_pr__nfet_01v8_59MFY5  sky130_fd_pr__nfet_01v8_59MFY5_2
timestamp 1641609411
transform 1 0 -91 0 1 -199
box -99 -157 99 157
use sky130_fd_pr__nfet_01v8_59MFY5  sky130_fd_pr__nfet_01v8_59MFY5_3
timestamp 1641609411
transform 1 0 -291 0 1 -199
box -99 -157 99 157
use sky130_fd_pr__pfet_01v8_MA8JHN  sky130_fd_pr__pfet_01v8_MA8JHN_0
timestamp 1641609411
transform 1 0 909 0 1 198
box -109 -198 109 164
use sky130_fd_pr__pfet_01v8_MA8JHN  sky130_fd_pr__pfet_01v8_MA8JHN_1
timestamp 1641609411
transform 1 0 709 0 1 198
box -109 -198 109 164
use sky130_fd_pr__pfet_01v8_MA8JHN  sky130_fd_pr__pfet_01v8_MA8JHN_2
timestamp 1641609411
transform 1 0 309 0 1 198
box -109 -198 109 164
use sky130_fd_pr__pfet_01v8_MA8JHN  sky130_fd_pr__pfet_01v8_MA8JHN_3
timestamp 1641609411
transform 1 0 109 0 1 198
box -109 -198 109 164
use sky130_fd_pr__pfet_01v8_MA8JHN  sky130_fd_pr__pfet_01v8_MA8JHN_4
timestamp 1641609411
transform 1 0 -491 0 1 198
box -109 -198 109 164
use sky130_fd_pr__pfet_01v8_MA8JHN  sky130_fd_pr__pfet_01v8_MA8JHN_5
timestamp 1641609411
transform 1 0 -291 0 1 198
box -109 -198 109 164
<< labels >>
flabel metal2 s 208 506 208 506 0 FreeSans 600 0 0 0 VDD
port 1 nsew
flabel metal1 s 216 -542 216 -542 0 FreeSans 600 0 0 0 GND
port 2 nsew
flabel metal2 s -284 -436 -284 -436 0 FreeSans 600 0 0 0 CLK
port 3 nsew
flabel metal1 s 904 328 904 328 0 FreeSans 600 0 0 0 IN
port 4 nsew
flabel metal1 s 8 320 8 320 0 FreeSans 600 0 0 0 ND
port 5 nsew
flabel locali s 400 320 400 320 0 FreeSans 600 0 0 0 D
port 6 nsew
<< end >>
