magic
tech sky130A
magscale 1 2
timestamp 1640975112
<< error_p >>
rect -28 144 28 150
rect -32 110 32 144
rect -28 104 28 110
rect 14 -162 16 94
<< nwell >>
rect -108 -198 108 164
<< pmos >>
rect -14 -136 14 64
<< pdiff >>
rect -72 49 -14 64
rect -72 15 -60 49
rect -26 15 -14 49
rect -72 -19 -14 15
rect -72 -53 -60 -19
rect -26 -53 -14 -19
rect -72 -87 -14 -53
rect -72 -121 -60 -87
rect -26 -121 -14 -87
rect -72 -136 -14 -121
rect 14 49 72 64
rect 14 15 26 49
rect 60 15 72 49
rect 14 -19 72 15
rect 14 -53 26 -19
rect 60 -53 72 -19
rect 14 -87 72 -53
rect 14 -121 26 -87
rect 60 -121 72 -87
rect 14 -136 72 -121
<< pdiffc >>
rect -60 15 -26 49
rect -60 -53 -26 -19
rect -60 -121 -26 -87
rect 26 15 60 49
rect 26 -53 60 -19
rect 26 -121 60 -87
<< poly >>
rect -32 94 32 160
rect -14 64 14 94
rect -14 -162 14 -136
<< locali >>
rect -32 110 32 144
rect -60 49 -26 68
rect -60 -19 -26 -17
rect -60 -55 -26 -53
rect -60 -140 -26 -121
rect 26 49 60 68
rect 26 -19 60 -17
rect 26 -55 60 -53
rect 26 -140 60 -121
<< viali >>
rect -60 15 -26 17
rect -60 -17 -26 15
rect -60 -87 -26 -55
rect -60 -89 -26 -87
rect 26 15 60 17
rect 26 -17 60 15
rect 26 -87 60 -55
rect 26 -89 60 -87
<< metal1 >>
rect -28 104 28 150
rect -66 17 -20 64
rect -66 -17 -60 17
rect -26 -17 -20 17
rect -66 -55 -20 -17
rect -66 -89 -60 -55
rect -26 -89 -20 -55
rect -66 -136 -20 -89
rect 20 17 66 64
rect 20 -17 26 17
rect 60 -17 66 17
rect 20 -55 66 -17
rect 20 -89 26 -55
rect 60 -89 66 -55
rect 20 -136 66 -89
<< end >>
