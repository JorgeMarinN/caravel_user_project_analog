magic
tech sky130A
magscale 1 2
timestamp 1640975112
<< nwell >>
rect -300 250 170 530
<< pwell >>
rect -286 -46 156 206
<< nmos >>
rect -20 -20 10 180
<< pmos >>
rect -20 290 10 490
<< ndiff >>
rect -140 131 -20 180
rect -140 97 -97 131
rect -63 97 -20 131
rect -140 63 -20 97
rect -140 29 -97 63
rect -63 29 -20 63
rect -140 -20 -20 29
rect 10 131 130 180
rect 10 97 53 131
rect 87 97 130 131
rect 10 63 130 97
rect 10 29 53 63
rect 87 29 130 63
rect 10 -20 130 29
<< pdiff >>
rect -140 441 -20 490
rect -140 407 -97 441
rect -63 407 -20 441
rect -140 373 -20 407
rect -140 339 -97 373
rect -63 339 -20 373
rect -140 290 -20 339
rect 10 441 130 490
rect 10 407 53 441
rect 87 407 130 441
rect 10 373 130 407
rect 10 339 53 373
rect 87 339 130 373
rect 10 290 130 339
<< ndiffc >>
rect -97 97 -63 131
rect -97 29 -63 63
rect 53 97 87 131
rect 53 29 87 63
<< pdiffc >>
rect -97 407 -63 441
rect -97 339 -63 373
rect 53 407 87 441
rect 53 339 87 373
<< psubdiff >>
rect -260 131 -140 180
rect -260 97 -217 131
rect -183 97 -140 131
rect -260 63 -140 97
rect -260 29 -217 63
rect -183 29 -140 63
rect -260 -20 -140 29
<< nsubdiff >>
rect -260 441 -140 490
rect -260 407 -217 441
rect -183 407 -140 441
rect -260 373 -140 407
rect -260 339 -217 373
rect -183 339 -140 373
rect -260 290 -140 339
<< psubdiffcont >>
rect -217 97 -183 131
rect -217 29 -183 63
<< nsubdiffcont >>
rect -217 407 -183 441
rect -217 339 -183 373
<< poly >>
rect -20 490 10 520
rect -20 180 10 290
rect -20 -50 10 -20
rect -90 -83 10 -50
rect -90 -117 -57 -83
rect -23 -117 10 -83
rect -90 -150 10 -117
<< polycont >>
rect -57 -117 -23 -83
<< locali >>
rect -250 443 -30 480
rect -250 407 -217 443
rect -183 407 -97 443
rect -63 407 -30 443
rect -250 373 -30 407
rect -250 337 -217 373
rect -183 337 -97 373
rect -63 337 -30 373
rect -250 300 -30 337
rect 20 441 120 480
rect 20 407 53 441
rect 87 407 120 441
rect 20 373 120 407
rect 20 339 53 373
rect 87 339 120 373
rect 20 300 120 339
rect 70 170 120 300
rect -250 133 -30 170
rect -250 97 -217 133
rect -183 97 -97 133
rect -63 97 -30 133
rect -250 63 -30 97
rect -250 27 -217 63
rect -183 27 -97 63
rect -63 27 -30 63
rect -250 -10 -30 27
rect 20 131 120 170
rect 20 97 53 131
rect 87 97 120 131
rect 20 63 120 97
rect 20 29 53 63
rect 87 29 120 63
rect 20 -10 120 29
rect 70 -50 120 -10
rect -300 -83 10 -50
rect -300 -100 -57 -83
rect -90 -117 -57 -100
rect -23 -117 10 -83
rect 70 -100 170 -50
rect -90 -150 10 -117
<< viali >>
rect -217 441 -183 443
rect -217 409 -183 441
rect -97 441 -63 443
rect -97 409 -63 441
rect -217 339 -183 371
rect -217 337 -183 339
rect -97 339 -63 371
rect -97 337 -63 339
rect -217 131 -183 133
rect -217 99 -183 131
rect -97 131 -63 133
rect -97 99 -63 131
rect -217 29 -183 61
rect -217 27 -183 29
rect -97 29 -63 61
rect -97 27 -63 29
<< metal1 >>
rect -300 443 170 480
rect -300 409 -217 443
rect -183 409 -97 443
rect -63 409 170 443
rect -300 371 170 409
rect -300 337 -217 371
rect -183 337 -97 371
rect -63 337 170 371
rect -300 300 170 337
rect -300 133 170 170
rect -300 99 -217 133
rect -183 99 -97 133
rect -63 99 170 133
rect -300 61 170 99
rect -300 27 -217 61
rect -183 27 -97 61
rect -63 27 170 61
rect -300 -10 170 27
<< labels >>
rlabel locali s -300 -80 -300 -80 4 VIN
port 1 nsew
rlabel locali s 170 -80 170 -80 4 VOUT
port 2 nsew
rlabel metal1 s -300 390 -300 390 4 VDD
port 3 nsew
rlabel metal1 s -300 80 -300 80 4 VSS
port 4 nsew
<< end >>
