magic
tech sky130A
magscale 1 2
timestamp 1641611256
<< nwell >>
rect -636 294 982 904
<< pwell >>
rect -472 -204 818 -70
<< psubdiff >>
rect -446 -120 792 -96
rect -446 -154 -422 -120
rect -388 -154 -354 -120
rect -320 -154 -286 -120
rect -252 -154 -218 -120
rect -184 -154 -150 -120
rect -116 -154 -82 -120
rect -48 -154 -14 -120
rect 20 -154 54 -120
rect 88 -154 122 -120
rect 156 -154 190 -120
rect 224 -154 258 -120
rect 292 -154 326 -120
rect 360 -154 394 -120
rect 428 -154 462 -120
rect 496 -154 530 -120
rect 564 -154 598 -120
rect 632 -154 666 -120
rect 700 -154 734 -120
rect 768 -154 792 -120
rect -446 -178 792 -154
<< nsubdiff >>
rect 2 824 336 852
rect 2 790 50 824
rect 84 790 118 824
rect 152 790 186 824
rect 220 790 254 824
rect 288 790 336 824
rect 2 692 336 790
<< psubdiffcont >>
rect -422 -154 -388 -120
rect -354 -154 -320 -120
rect -286 -154 -252 -120
rect -218 -154 -184 -120
rect -150 -154 -116 -120
rect -82 -154 -48 -120
rect -14 -154 20 -120
rect 54 -154 88 -120
rect 122 -154 156 -120
rect 190 -154 224 -120
rect 258 -154 292 -120
rect 326 -154 360 -120
rect 394 -154 428 -120
rect 462 -154 496 -120
rect 530 -154 564 -120
rect 598 -154 632 -120
rect 666 -154 700 -120
rect 734 -154 768 -120
<< nsubdiffcont >>
rect 50 790 84 824
rect 118 790 152 824
rect 186 790 220 824
rect 254 790 288 824
<< poly >>
rect -542 226 -512 356
rect 58 252 88 330
rect 258 252 288 330
rect 858 226 888 356
<< locali >>
rect 14 824 324 840
rect 14 790 44 824
rect 84 790 116 824
rect 152 790 186 824
rect 222 790 254 824
rect 294 790 324 824
rect 14 774 324 790
rect 50 692 400 738
rect -678 602 -494 638
rect 50 604 96 692
rect -678 316 -644 602
rect 354 560 400 692
rect 334 522 400 560
rect 612 316 646 352
rect -678 282 646 316
rect -440 -120 786 -96
rect -440 -154 -422 -120
rect -386 -154 -354 -120
rect -314 -154 -286 -120
rect -242 -154 -218 -120
rect -170 -154 -150 -120
rect -98 -154 -82 -120
rect -26 -154 -14 -120
rect 46 -154 54 -120
rect 118 -154 122 -120
rect 224 -154 228 -120
rect 292 -154 300 -120
rect 360 -154 372 -120
rect 428 -154 444 -120
rect 496 -154 516 -120
rect 564 -154 588 -120
rect 632 -154 660 -120
rect 700 -154 732 -120
rect 768 -154 786 -120
rect -440 -174 786 -154
<< viali >>
rect 44 790 50 824
rect 50 790 78 824
rect 116 790 118 824
rect 118 790 150 824
rect 188 790 220 824
rect 220 790 222 824
rect 260 790 288 824
rect 288 790 294 824
rect -420 -154 -388 -120
rect -388 -154 -386 -120
rect -348 -154 -320 -120
rect -320 -154 -314 -120
rect -276 -154 -252 -120
rect -252 -154 -242 -120
rect -204 -154 -184 -120
rect -184 -154 -170 -120
rect -132 -154 -116 -120
rect -116 -154 -98 -120
rect -60 -154 -48 -120
rect -48 -154 -26 -120
rect 12 -154 20 -120
rect 20 -154 46 -120
rect 84 -154 88 -120
rect 88 -154 118 -120
rect 156 -154 190 -120
rect 228 -154 258 -120
rect 258 -154 262 -120
rect 300 -154 326 -120
rect 326 -154 334 -120
rect 372 -154 394 -120
rect 394 -154 406 -120
rect 444 -154 462 -120
rect 462 -154 478 -120
rect 516 -154 530 -120
rect 530 -154 550 -120
rect 588 -154 598 -120
rect 598 -154 622 -120
rect 660 -154 666 -120
rect 666 -154 694 -120
rect 732 -154 734 -120
rect 734 -154 766 -120
<< metal1 >>
rect 138 842 208 848
rect 138 840 147 842
rect -640 824 147 840
rect 199 840 208 842
rect 199 824 986 840
rect -640 790 44 824
rect 78 790 116 824
rect 222 790 260 824
rect 294 790 986 824
rect -640 776 986 790
rect -640 356 -594 776
rect 14 774 324 776
rect -60 692 296 738
rect -550 655 -486 662
rect -550 654 -544 655
rect -560 603 -544 654
rect -492 603 -486 655
rect -350 655 -286 662
rect -350 654 -344 655
rect -560 596 -486 603
rect -360 603 -344 654
rect -292 603 -286 655
rect -360 596 -286 603
rect -560 586 -494 596
rect -360 586 -294 596
rect -60 556 -14 692
rect 40 588 106 654
rect 250 652 296 692
rect 632 655 696 662
rect 240 586 306 652
rect 632 603 638 655
rect 690 654 696 655
rect 832 654 896 660
rect 690 603 706 654
rect 632 596 706 603
rect 832 602 838 654
rect 890 602 906 654
rect 832 596 906 602
rect 640 586 706 596
rect 840 586 906 596
rect -460 356 -394 556
rect -60 518 6 556
rect 140 541 206 556
rect 140 489 147 541
rect 199 489 206 541
rect 140 356 206 489
rect 740 356 806 556
rect 940 356 986 776
rect -600 316 -536 322
rect -306 316 -260 356
rect -600 264 -594 316
rect -542 266 -260 316
rect -542 264 -536 266
rect -600 258 -536 264
rect -594 226 -548 258
rect 6 226 52 356
rect 294 226 340 356
rect 606 316 652 356
rect 882 316 946 322
rect 606 266 888 316
rect 882 264 888 266
rect 940 264 946 316
rect 882 258 946 264
rect 894 226 940 258
rect -466 26 -394 226
rect -260 26 -194 226
rect -60 26 6 226
rect 140 26 206 226
rect 340 26 406 226
rect 540 26 606 226
rect 740 26 812 226
rect -440 -108 -394 26
rect -360 -6 -294 -4
rect -160 -6 -94 -4
rect -360 -12 -286 -6
rect -360 -62 -344 -12
rect -350 -64 -344 -62
rect -292 -64 -286 -12
rect -160 -12 -86 -6
rect -160 -62 -144 -12
rect -350 -70 -286 -64
rect -150 -64 -144 -62
rect -92 -64 -86 -12
rect -150 -70 -86 -64
rect 94 -108 252 26
rect 440 -6 506 -4
rect 640 -6 706 -4
rect 432 -12 506 -6
rect 432 -64 438 -12
rect 490 -62 506 -12
rect 632 -12 706 -6
rect 490 -64 496 -62
rect 432 -70 496 -64
rect 632 -64 638 -12
rect 690 -62 706 -12
rect 690 -64 696 -62
rect 632 -70 696 -64
rect 740 -108 786 26
rect -440 -120 786 -108
rect -440 -154 -420 -120
rect -386 -154 -348 -120
rect -314 -154 -276 -120
rect -242 -154 -204 -120
rect -170 -154 -132 -120
rect -98 -154 -60 -120
rect -26 -154 12 -120
rect 46 -154 84 -120
rect 118 -154 156 -120
rect 190 -154 228 -120
rect 262 -154 300 -120
rect 334 -154 372 -120
rect 406 -154 444 -120
rect 478 -154 516 -120
rect 550 -154 588 -120
rect 622 -154 660 -120
rect 694 -154 732 -120
rect 766 -154 786 -120
rect -440 -166 786 -154
<< via1 >>
rect 147 824 199 842
rect 147 790 150 824
rect 150 790 188 824
rect 188 790 199 824
rect -544 603 -492 655
rect -344 603 -292 655
rect 638 603 690 655
rect 838 602 890 654
rect 147 489 199 541
rect -594 264 -542 316
rect 888 264 940 316
rect -344 -64 -292 -12
rect -144 -64 -92 -12
rect 438 -64 490 -12
rect 638 -64 690 -12
<< metal2 >>
rect 138 842 208 848
rect 138 790 147 842
rect 199 790 208 842
rect 138 784 208 790
rect -550 655 -486 662
rect -550 603 -544 655
rect -492 603 -486 655
rect -550 596 -486 603
rect -350 655 -286 662
rect -350 603 -344 655
rect -292 603 -286 655
rect -350 440 -286 603
rect 150 548 196 784
rect 632 655 696 662
rect 632 603 638 655
rect 690 603 696 655
rect 140 541 206 548
rect 140 489 147 541
rect 199 489 206 541
rect 140 482 206 489
rect 632 440 696 603
rect 832 654 896 660
rect 832 602 838 654
rect 890 602 896 654
rect 832 596 896 602
rect -350 374 696 440
rect -600 316 -536 324
rect -600 264 -594 316
rect -542 264 -536 316
rect -600 -106 -536 264
rect 150 108 196 374
rect 882 316 946 322
rect 882 264 888 316
rect 940 264 946 316
rect -350 44 696 108
rect -350 -12 -286 44
rect -350 -64 -344 -12
rect -292 -64 -286 -12
rect -350 -70 -286 -64
rect -150 -12 -84 -6
rect -150 -64 -144 -12
rect -92 -64 -84 -12
rect -150 -106 -84 -64
rect -600 -166 -84 -106
rect 432 -12 496 -6
rect 432 -64 438 -12
rect 490 -64 496 -12
rect 432 -106 496 -64
rect 632 -12 696 44
rect 632 -64 638 -12
rect 690 -64 696 -12
rect 632 -70 696 -64
rect 882 -106 946 264
rect 432 -166 946 -106
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_0
timestamp 1641609411
transform 1 0 -527 0 1 126
box -99 -126 99 126
use sky130_fd_pr__pfet_01v8_MA8JHN  sky130_fd_pr__pfet_01v8_MA8JHN_1
timestamp 1641609411
transform 1 0 -527 0 1 492
box -109 -198 109 164
use sky130_fd_pr__pfet_01v8_MA8JHN  sky130_fd_pr__pfet_01v8_MA8JHN_0
timestamp 1641609411
transform 1 0 -327 0 1 492
box -109 -198 109 164
use sky130_fd_pr__nfet_01v8_59MFY5  sky130_fd_pr__nfet_01v8_59MFY5_0
timestamp 1641609411
transform 1 0 -327 0 1 95
box -99 -157 99 157
use sky130_fd_pr__nfet_01v8_59MFY5  sky130_fd_pr__nfet_01v8_59MFY5_1
timestamp 1641609411
transform 1 0 -127 0 1 95
box -99 -157 99 157
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_1
timestamp 1641609411
transform 1 0 73 0 1 126
box -99 -126 99 126
use sky130_fd_pr__pfet_01v8_MA8JHN  sky130_fd_pr__pfet_01v8_MA8JHN_2
timestamp 1641609411
transform 1 0 73 0 1 492
box -109 -198 109 164
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_2
timestamp 1641609411
transform 1 0 273 0 1 126
box -99 -126 99 126
use sky130_fd_pr__pfet_01v8_MA8JHN  sky130_fd_pr__pfet_01v8_MA8JHN_3
timestamp 1641609411
transform 1 0 273 0 1 492
box -109 -198 109 164
use sky130_fd_pr__nfet_01v8_59MFY5  sky130_fd_pr__nfet_01v8_59MFY5_2
timestamp 1641609411
transform 1 0 473 0 1 95
box -99 -157 99 157
use sky130_fd_pr__pfet_01v8_MA8JHN  sky130_fd_pr__pfet_01v8_MA8JHN_4
timestamp 1641609411
transform 1 0 673 0 1 492
box -109 -198 109 164
use sky130_fd_pr__nfet_01v8_59MFY5  sky130_fd_pr__nfet_01v8_59MFY5_3
timestamp 1641609411
transform 1 0 673 0 1 95
box -99 -157 99 157
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_3
timestamp 1641609411
transform 1 0 873 0 1 126
box -99 -126 99 126
use sky130_fd_pr__pfet_01v8_MA8JHN  sky130_fd_pr__pfet_01v8_MA8JHN_5
timestamp 1641609411
transform 1 0 873 0 1 492
box -109 -198 109 164
<< labels >>
flabel metal2 s 476 -40 476 -40 0 FreeSans 600 0 0 0 NDIFF
port 1 nsew
flabel metal2 s -120 -32 -120 -32 0 FreeSans 600 0 0 0 PDIFF
port 2 nsew
flabel metal2 s 172 758 172 758 0 FreeSans 600 0 0 0 VDD
port 3 nsew
flabel metal2 s 170 76 170 76 0 FreeSans 600 0 0 0 CLK
port 4 nsew
flabel metal1 s -40 630 -40 630 0 FreeSans 600 0 0 0 ND
port 5 nsew
flabel locali s 380 624 380 624 0 FreeSans 600 0 0 0 D
port 6 nsew
flabel metal1 s 168 -76 168 -76 0 FreeSans 600 0 0 0 GND
port 7 nsew
flabel metal2 s 868 624 868 624 0 FreeSans 600 0 0 0 IN
port 8 nsew
<< end >>
