magic
tech sky130A
magscale 1 2
timestamp 1641609411
<< metal4 >>
rect -671 2198 671 2320
rect -671 1962 415 2198
rect 651 1962 671 2198
rect -671 1878 671 1962
rect -671 1642 415 1878
rect 651 1642 671 1878
rect -671 1558 671 1642
rect -671 1322 415 1558
rect 651 1322 671 1558
rect -671 1238 671 1322
rect -671 1002 415 1238
rect 651 1002 671 1238
rect -671 918 671 1002
rect -671 682 415 918
rect 651 682 671 918
rect -671 598 671 682
rect -671 362 415 598
rect 651 362 671 598
rect -671 278 671 362
rect -671 42 415 278
rect 651 42 671 278
rect -671 -42 671 42
rect -671 -278 415 -42
rect 651 -278 671 -42
rect -671 -362 671 -278
rect -671 -598 415 -362
rect 651 -598 671 -362
rect -671 -682 671 -598
rect -671 -918 415 -682
rect 651 -918 671 -682
rect -671 -1002 671 -918
rect -671 -1238 415 -1002
rect 651 -1238 671 -1002
rect -671 -1322 671 -1238
rect -671 -1558 415 -1322
rect 651 -1558 671 -1322
rect -671 -1642 671 -1558
rect -671 -1878 415 -1642
rect 651 -1878 671 -1642
rect -671 -1962 671 -1878
rect -671 -2198 415 -1962
rect 651 -2198 671 -1962
rect -671 -2320 671 -2198
<< via4 >>
rect 415 1962 651 2198
rect 415 1642 651 1878
rect 415 1322 651 1558
rect 415 1002 651 1238
rect 415 682 651 918
rect 415 362 651 598
rect 415 42 651 278
rect 415 -278 651 -42
rect 415 -598 651 -362
rect 415 -918 651 -682
rect 415 -1238 651 -1002
rect 415 -1558 651 -1322
rect 415 -1878 651 -1642
rect 415 -2198 651 -1962
<< mimcap2 >>
rect -571 2038 69 2220
rect -571 -2038 -529 2038
rect 27 -2038 69 2038
rect -571 -2220 69 -2038
<< mimcap2contact >>
rect -529 -2038 27 2038
<< metal5 >>
rect -555 2038 53 2204
rect -555 -2038 -529 2038
rect 27 -2038 53 2038
rect -555 -2204 53 -2038
rect 373 2198 693 2321
rect 373 1962 415 2198
rect 651 1962 693 2198
rect 373 1878 693 1962
rect 373 1642 415 1878
rect 651 1642 693 1878
rect 373 1558 693 1642
rect 373 1322 415 1558
rect 651 1322 693 1558
rect 373 1238 693 1322
rect 373 1002 415 1238
rect 651 1002 693 1238
rect 373 918 693 1002
rect 373 682 415 918
rect 651 682 693 918
rect 373 598 693 682
rect 373 362 415 598
rect 651 362 693 598
rect 373 278 693 362
rect 373 42 415 278
rect 651 42 693 278
rect 373 -42 693 42
rect 373 -278 415 -42
rect 651 -278 693 -42
rect 373 -362 693 -278
rect 373 -598 415 -362
rect 651 -598 693 -362
rect 373 -682 693 -598
rect 373 -918 415 -682
rect 651 -918 693 -682
rect 373 -1002 693 -918
rect 373 -1238 415 -1002
rect 651 -1238 693 -1002
rect 373 -1322 693 -1238
rect 373 -1558 415 -1322
rect 651 -1558 693 -1322
rect 373 -1642 693 -1558
rect 373 -1878 415 -1642
rect 651 -1878 693 -1642
rect 373 -1962 693 -1878
rect 373 -2198 415 -1962
rect 651 -2198 693 -1962
rect 373 -2321 693 -2198
<< properties >>
string FIXED_BBOX -671 -2320 169 2320
<< end >>
