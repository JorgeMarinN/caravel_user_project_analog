magic
tech sky130A
magscale 1 2
timestamp 1641609411
<< metal3 >>
rect -456 2272 456 2320
rect -456 2208 372 2272
rect 436 2208 456 2272
rect -456 2192 456 2208
rect -456 2128 372 2192
rect 436 2128 456 2192
rect -456 2112 456 2128
rect -456 2048 372 2112
rect 436 2048 456 2112
rect -456 2032 456 2048
rect -456 1968 372 2032
rect 436 1968 456 2032
rect -456 1952 456 1968
rect -456 1888 372 1952
rect 436 1888 456 1952
rect -456 1872 456 1888
rect -456 1808 372 1872
rect 436 1808 456 1872
rect -456 1792 456 1808
rect -456 1728 372 1792
rect 436 1728 456 1792
rect -456 1712 456 1728
rect -456 1648 372 1712
rect 436 1648 456 1712
rect -456 1632 456 1648
rect -456 1568 372 1632
rect 436 1568 456 1632
rect -456 1552 456 1568
rect -456 1488 372 1552
rect 436 1488 456 1552
rect -456 1472 456 1488
rect -456 1408 372 1472
rect 436 1408 456 1472
rect -456 1392 456 1408
rect -456 1328 372 1392
rect 436 1328 456 1392
rect -456 1312 456 1328
rect -456 1248 372 1312
rect 436 1248 456 1312
rect -456 1232 456 1248
rect -456 1168 372 1232
rect 436 1168 456 1232
rect -456 1152 456 1168
rect -456 1088 372 1152
rect 436 1088 456 1152
rect -456 1072 456 1088
rect -456 1008 372 1072
rect 436 1008 456 1072
rect -456 992 456 1008
rect -456 928 372 992
rect 436 928 456 992
rect -456 912 456 928
rect -456 848 372 912
rect 436 848 456 912
rect -456 832 456 848
rect -456 768 372 832
rect 436 768 456 832
rect -456 752 456 768
rect -456 688 372 752
rect 436 688 456 752
rect -456 672 456 688
rect -456 608 372 672
rect 436 608 456 672
rect -456 592 456 608
rect -456 528 372 592
rect 436 528 456 592
rect -456 512 456 528
rect -456 448 372 512
rect 436 448 456 512
rect -456 432 456 448
rect -456 368 372 432
rect 436 368 456 432
rect -456 352 456 368
rect -456 288 372 352
rect 436 288 456 352
rect -456 272 456 288
rect -456 208 372 272
rect 436 208 456 272
rect -456 192 456 208
rect -456 128 372 192
rect 436 128 456 192
rect -456 112 456 128
rect -456 48 372 112
rect 436 48 456 112
rect -456 32 456 48
rect -456 -32 372 32
rect 436 -32 456 32
rect -456 -48 456 -32
rect -456 -112 372 -48
rect 436 -112 456 -48
rect -456 -128 456 -112
rect -456 -192 372 -128
rect 436 -192 456 -128
rect -456 -208 456 -192
rect -456 -272 372 -208
rect 436 -272 456 -208
rect -456 -288 456 -272
rect -456 -352 372 -288
rect 436 -352 456 -288
rect -456 -368 456 -352
rect -456 -432 372 -368
rect 436 -432 456 -368
rect -456 -448 456 -432
rect -456 -512 372 -448
rect 436 -512 456 -448
rect -456 -528 456 -512
rect -456 -592 372 -528
rect 436 -592 456 -528
rect -456 -608 456 -592
rect -456 -672 372 -608
rect 436 -672 456 -608
rect -456 -688 456 -672
rect -456 -752 372 -688
rect 436 -752 456 -688
rect -456 -768 456 -752
rect -456 -832 372 -768
rect 436 -832 456 -768
rect -456 -848 456 -832
rect -456 -912 372 -848
rect 436 -912 456 -848
rect -456 -928 456 -912
rect -456 -992 372 -928
rect 436 -992 456 -928
rect -456 -1008 456 -992
rect -456 -1072 372 -1008
rect 436 -1072 456 -1008
rect -456 -1088 456 -1072
rect -456 -1152 372 -1088
rect 436 -1152 456 -1088
rect -456 -1168 456 -1152
rect -456 -1232 372 -1168
rect 436 -1232 456 -1168
rect -456 -1248 456 -1232
rect -456 -1312 372 -1248
rect 436 -1312 456 -1248
rect -456 -1328 456 -1312
rect -456 -1392 372 -1328
rect 436 -1392 456 -1328
rect -456 -1408 456 -1392
rect -456 -1472 372 -1408
rect 436 -1472 456 -1408
rect -456 -1488 456 -1472
rect -456 -1552 372 -1488
rect 436 -1552 456 -1488
rect -456 -1568 456 -1552
rect -456 -1632 372 -1568
rect 436 -1632 456 -1568
rect -456 -1648 456 -1632
rect -456 -1712 372 -1648
rect 436 -1712 456 -1648
rect -456 -1728 456 -1712
rect -456 -1792 372 -1728
rect 436 -1792 456 -1728
rect -456 -1808 456 -1792
rect -456 -1872 372 -1808
rect 436 -1872 456 -1808
rect -456 -1888 456 -1872
rect -456 -1952 372 -1888
rect 436 -1952 456 -1888
rect -456 -1968 456 -1952
rect -456 -2032 372 -1968
rect 436 -2032 456 -1968
rect -456 -2048 456 -2032
rect -456 -2112 372 -2048
rect 436 -2112 456 -2048
rect -456 -2128 456 -2112
rect -456 -2192 372 -2128
rect 436 -2192 456 -2128
rect -456 -2208 456 -2192
rect -456 -2272 372 -2208
rect 436 -2272 456 -2208
rect -456 -2320 456 -2272
<< via3 >>
rect 372 2208 436 2272
rect 372 2128 436 2192
rect 372 2048 436 2112
rect 372 1968 436 2032
rect 372 1888 436 1952
rect 372 1808 436 1872
rect 372 1728 436 1792
rect 372 1648 436 1712
rect 372 1568 436 1632
rect 372 1488 436 1552
rect 372 1408 436 1472
rect 372 1328 436 1392
rect 372 1248 436 1312
rect 372 1168 436 1232
rect 372 1088 436 1152
rect 372 1008 436 1072
rect 372 928 436 992
rect 372 848 436 912
rect 372 768 436 832
rect 372 688 436 752
rect 372 608 436 672
rect 372 528 436 592
rect 372 448 436 512
rect 372 368 436 432
rect 372 288 436 352
rect 372 208 436 272
rect 372 128 436 192
rect 372 48 436 112
rect 372 -32 436 32
rect 372 -112 436 -48
rect 372 -192 436 -128
rect 372 -272 436 -208
rect 372 -352 436 -288
rect 372 -432 436 -368
rect 372 -512 436 -448
rect 372 -592 436 -528
rect 372 -672 436 -608
rect 372 -752 436 -688
rect 372 -832 436 -768
rect 372 -912 436 -848
rect 372 -992 436 -928
rect 372 -1072 436 -1008
rect 372 -1152 436 -1088
rect 372 -1232 436 -1168
rect 372 -1312 436 -1248
rect 372 -1392 436 -1328
rect 372 -1472 436 -1408
rect 372 -1552 436 -1488
rect 372 -1632 436 -1568
rect 372 -1712 436 -1648
rect 372 -1792 436 -1728
rect 372 -1872 436 -1808
rect 372 -1952 436 -1888
rect 372 -2032 436 -1968
rect 372 -2112 436 -2048
rect 372 -2192 436 -2128
rect 372 -2272 436 -2208
<< mimcap >>
rect -356 2152 284 2220
rect -356 -2152 -68 2152
rect -4 -2152 284 2152
rect -356 -2220 284 -2152
<< mimcapcontact >>
rect -68 -2152 -4 2152
<< metal4 >>
rect 356 2272 452 2308
rect 356 2208 372 2272
rect 436 2208 452 2272
rect 356 2192 452 2208
rect -69 2152 -3 2181
rect -69 -2152 -68 2152
rect -4 -2152 -3 2152
rect -69 -2181 -3 -2152
rect 356 2128 372 2192
rect 436 2128 452 2192
rect 356 2112 452 2128
rect 356 2048 372 2112
rect 436 2048 452 2112
rect 356 2032 452 2048
rect 356 1968 372 2032
rect 436 1968 452 2032
rect 356 1952 452 1968
rect 356 1888 372 1952
rect 436 1888 452 1952
rect 356 1872 452 1888
rect 356 1808 372 1872
rect 436 1808 452 1872
rect 356 1792 452 1808
rect 356 1728 372 1792
rect 436 1728 452 1792
rect 356 1712 452 1728
rect 356 1648 372 1712
rect 436 1648 452 1712
rect 356 1632 452 1648
rect 356 1568 372 1632
rect 436 1568 452 1632
rect 356 1552 452 1568
rect 356 1488 372 1552
rect 436 1488 452 1552
rect 356 1472 452 1488
rect 356 1408 372 1472
rect 436 1408 452 1472
rect 356 1392 452 1408
rect 356 1328 372 1392
rect 436 1328 452 1392
rect 356 1312 452 1328
rect 356 1248 372 1312
rect 436 1248 452 1312
rect 356 1232 452 1248
rect 356 1168 372 1232
rect 436 1168 452 1232
rect 356 1152 452 1168
rect 356 1088 372 1152
rect 436 1088 452 1152
rect 356 1072 452 1088
rect 356 1008 372 1072
rect 436 1008 452 1072
rect 356 992 452 1008
rect 356 928 372 992
rect 436 928 452 992
rect 356 912 452 928
rect 356 848 372 912
rect 436 848 452 912
rect 356 832 452 848
rect 356 768 372 832
rect 436 768 452 832
rect 356 752 452 768
rect 356 688 372 752
rect 436 688 452 752
rect 356 672 452 688
rect 356 608 372 672
rect 436 608 452 672
rect 356 592 452 608
rect 356 528 372 592
rect 436 528 452 592
rect 356 512 452 528
rect 356 448 372 512
rect 436 448 452 512
rect 356 432 452 448
rect 356 368 372 432
rect 436 368 452 432
rect 356 352 452 368
rect 356 288 372 352
rect 436 288 452 352
rect 356 272 452 288
rect 356 208 372 272
rect 436 208 452 272
rect 356 192 452 208
rect 356 128 372 192
rect 436 128 452 192
rect 356 112 452 128
rect 356 48 372 112
rect 436 48 452 112
rect 356 32 452 48
rect 356 -32 372 32
rect 436 -32 452 32
rect 356 -48 452 -32
rect 356 -112 372 -48
rect 436 -112 452 -48
rect 356 -128 452 -112
rect 356 -192 372 -128
rect 436 -192 452 -128
rect 356 -208 452 -192
rect 356 -272 372 -208
rect 436 -272 452 -208
rect 356 -288 452 -272
rect 356 -352 372 -288
rect 436 -352 452 -288
rect 356 -368 452 -352
rect 356 -432 372 -368
rect 436 -432 452 -368
rect 356 -448 452 -432
rect 356 -512 372 -448
rect 436 -512 452 -448
rect 356 -528 452 -512
rect 356 -592 372 -528
rect 436 -592 452 -528
rect 356 -608 452 -592
rect 356 -672 372 -608
rect 436 -672 452 -608
rect 356 -688 452 -672
rect 356 -752 372 -688
rect 436 -752 452 -688
rect 356 -768 452 -752
rect 356 -832 372 -768
rect 436 -832 452 -768
rect 356 -848 452 -832
rect 356 -912 372 -848
rect 436 -912 452 -848
rect 356 -928 452 -912
rect 356 -992 372 -928
rect 436 -992 452 -928
rect 356 -1008 452 -992
rect 356 -1072 372 -1008
rect 436 -1072 452 -1008
rect 356 -1088 452 -1072
rect 356 -1152 372 -1088
rect 436 -1152 452 -1088
rect 356 -1168 452 -1152
rect 356 -1232 372 -1168
rect 436 -1232 452 -1168
rect 356 -1248 452 -1232
rect 356 -1312 372 -1248
rect 436 -1312 452 -1248
rect 356 -1328 452 -1312
rect 356 -1392 372 -1328
rect 436 -1392 452 -1328
rect 356 -1408 452 -1392
rect 356 -1472 372 -1408
rect 436 -1472 452 -1408
rect 356 -1488 452 -1472
rect 356 -1552 372 -1488
rect 436 -1552 452 -1488
rect 356 -1568 452 -1552
rect 356 -1632 372 -1568
rect 436 -1632 452 -1568
rect 356 -1648 452 -1632
rect 356 -1712 372 -1648
rect 436 -1712 452 -1648
rect 356 -1728 452 -1712
rect 356 -1792 372 -1728
rect 436 -1792 452 -1728
rect 356 -1808 452 -1792
rect 356 -1872 372 -1808
rect 436 -1872 452 -1808
rect 356 -1888 452 -1872
rect 356 -1952 372 -1888
rect 436 -1952 452 -1888
rect 356 -1968 452 -1952
rect 356 -2032 372 -1968
rect 436 -2032 452 -1968
rect 356 -2048 452 -2032
rect 356 -2112 372 -2048
rect 436 -2112 452 -2048
rect 356 -2128 452 -2112
rect 356 -2192 372 -2128
rect 436 -2192 452 -2128
rect 356 -2208 452 -2192
rect 356 -2272 372 -2208
rect 436 -2272 452 -2208
rect 356 -2308 452 -2272
<< properties >>
string FIXED_BBOX -456 -2320 384 2320
<< end >>
