magic
tech sky130A
magscale 1 2
timestamp 1641609411
<< error_p >>
rect -29 145 29 151
rect -29 111 -17 145
rect -29 105 29 111
<< nwell >>
rect -109 -198 109 164
<< pmos >>
rect -15 -136 15 64
<< pdiff >>
rect -73 49 -15 64
rect -73 15 -61 49
rect -27 15 -15 49
rect -73 -19 -15 15
rect -73 -53 -61 -19
rect -27 -53 -15 -19
rect -73 -87 -15 -53
rect -73 -121 -61 -87
rect -27 -121 -15 -87
rect -73 -136 -15 -121
rect 15 49 73 64
rect 15 15 27 49
rect 61 15 73 49
rect 15 -19 73 15
rect 15 -53 27 -19
rect 61 -53 73 -19
rect 15 -87 73 -53
rect 15 -121 27 -87
rect 61 -121 73 -87
rect 15 -136 73 -121
<< pdiffc >>
rect -61 15 -27 49
rect -61 -53 -27 -19
rect -61 -121 -27 -87
rect 27 15 61 49
rect 27 -53 61 -19
rect 27 -121 61 -87
<< poly >>
rect -33 145 33 161
rect -33 111 -17 145
rect 17 111 33 145
rect -33 95 33 111
rect -15 64 15 95
rect -15 -162 15 -136
<< polycont >>
rect -17 111 17 145
<< locali >>
rect -33 111 -17 145
rect 17 111 33 145
rect -61 49 -27 68
rect -61 -19 -27 -17
rect -61 -55 -27 -53
rect -61 -140 -27 -121
rect 27 49 61 68
rect 27 -19 61 -17
rect 27 -55 61 -53
rect 27 -140 61 -121
<< viali >>
rect -17 111 17 145
rect -61 15 -27 17
rect -61 -17 -27 15
rect -61 -87 -27 -55
rect -61 -89 -27 -87
rect 27 15 61 17
rect 27 -17 61 15
rect 27 -87 61 -55
rect 27 -89 61 -87
<< metal1 >>
rect -29 145 29 151
rect -29 111 -17 145
rect 17 111 29 145
rect -29 105 29 111
rect -67 17 -21 64
rect -67 -17 -61 17
rect -27 -17 -21 17
rect -67 -55 -21 -17
rect -67 -89 -61 -55
rect -27 -89 -21 -55
rect -67 -136 -21 -89
rect 21 17 67 64
rect 21 -17 27 17
rect 61 -17 67 17
rect 21 -55 67 -17
rect 21 -89 27 -55
rect 61 -89 67 -55
rect 21 -136 67 -89
<< end >>
