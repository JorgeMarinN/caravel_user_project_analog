magic
tech sky130A
magscale 1 2
timestamp 1640991954
<< metal2 >>
rect 9938 4588 10022 4622
rect 9938 4532 9952 4588
rect 10008 4532 10022 4588
rect 9938 4508 10022 4532
rect 9938 4452 9952 4508
rect 10008 4452 10022 4508
rect 9938 4428 10022 4452
rect 9938 4372 9952 4428
rect 10008 4372 10022 4428
rect 9938 4348 10022 4372
rect 9938 4292 9952 4348
rect 10008 4292 10022 4348
rect 9938 4268 10022 4292
rect 9938 4212 9952 4268
rect 10008 4212 10022 4268
rect 9938 4188 10022 4212
rect 9938 4132 9952 4188
rect 10008 4132 10022 4188
rect 9938 4108 10022 4132
rect 9938 4052 9952 4108
rect 10008 4052 10022 4108
rect 9938 4028 10022 4052
rect 9938 3972 9952 4028
rect 10008 3972 10022 4028
rect 9938 3948 10022 3972
rect 9938 3892 9952 3948
rect 10008 3892 10022 3948
rect 9938 3868 10022 3892
rect 9938 3812 9952 3868
rect 10008 3812 10022 3868
rect 9938 3788 10022 3812
rect 9938 3732 9952 3788
rect 10008 3732 10022 3788
rect 9938 3708 10022 3732
rect 9938 3652 9952 3708
rect 10008 3652 10022 3708
rect 9938 3628 10022 3652
rect 9938 3572 9952 3628
rect 10008 3572 10022 3628
rect 9938 3548 10022 3572
rect 9938 3492 9952 3548
rect 10008 3492 10022 3548
rect 9938 3468 10022 3492
rect 9938 3412 9952 3468
rect 10008 3412 10022 3468
rect 9938 3388 10022 3412
rect 9938 3332 9952 3388
rect 10008 3332 10022 3388
rect 9938 3308 10022 3332
rect 9938 3252 9952 3308
rect 10008 3252 10022 3308
rect 9938 3228 10022 3252
rect 9938 3172 9952 3228
rect 10008 3172 10022 3228
rect 9938 3148 10022 3172
rect 9938 3092 9952 3148
rect 10008 3092 10022 3148
rect 9938 3068 10022 3092
rect 9938 3012 9952 3068
rect 10008 3012 10022 3068
rect 9938 2988 10022 3012
rect 9938 2932 9952 2988
rect 10008 2932 10022 2988
rect 9938 2908 10022 2932
rect 9938 2852 9952 2908
rect 10008 2852 10022 2908
rect 9938 2828 10022 2852
rect 9938 2772 9952 2828
rect 10008 2772 10022 2828
rect 9938 2748 10022 2772
rect 9938 2692 9952 2748
rect 10008 2692 10022 2748
rect 9938 2668 10022 2692
rect 9938 2612 9952 2668
rect 10008 2612 10022 2668
rect 9938 2588 10022 2612
rect 9938 2532 9952 2588
rect 10008 2532 10022 2588
rect 9938 2508 10022 2532
rect 9938 2452 9952 2508
rect 10008 2452 10022 2508
rect 9938 2428 10022 2452
rect 9938 2372 9952 2428
rect 10008 2372 10022 2428
rect 9938 2348 10022 2372
rect 9938 2292 9952 2348
rect 10008 2292 10022 2348
rect 9938 2268 10022 2292
rect 9938 2212 9952 2268
rect 10008 2212 10022 2268
rect 9938 2188 10022 2212
rect 9938 2132 9952 2188
rect 10008 2132 10022 2188
rect 9938 2108 10022 2132
rect 9938 2052 9952 2108
rect 10008 2052 10022 2108
rect 9938 2028 10022 2052
rect 9938 1972 9952 2028
rect 10008 1972 10022 2028
rect 9938 1948 10022 1972
rect 9938 1892 9952 1948
rect 10008 1892 10022 1948
rect 9938 1868 10022 1892
rect 9938 1812 9952 1868
rect 10008 1812 10022 1868
rect 9938 1788 10022 1812
rect 9938 1732 9952 1788
rect 10008 1732 10022 1788
rect 9938 1708 10022 1732
rect 9938 1652 9952 1708
rect 10008 1652 10022 1708
rect 9938 1628 10022 1652
rect 9938 1572 9952 1628
rect 10008 1572 10022 1628
rect 9938 1548 10022 1572
rect 9938 1492 9952 1548
rect 10008 1492 10022 1548
rect 9938 1468 10022 1492
rect 9938 1412 9952 1468
rect 10008 1412 10022 1468
rect 9938 1388 10022 1412
rect 9938 1332 9952 1388
rect 10008 1332 10022 1388
rect 9938 1308 10022 1332
rect 9938 1252 9952 1308
rect 10008 1252 10022 1308
rect 9938 1228 10022 1252
rect 9938 1172 9952 1228
rect 10008 1172 10022 1228
rect 9938 1148 10022 1172
rect 9938 1092 9952 1148
rect 10008 1092 10022 1148
rect 9938 1068 10022 1092
rect 9938 1012 9952 1068
rect 10008 1012 10022 1068
rect 9938 988 10022 1012
rect 9938 932 9952 988
rect 10008 932 10022 988
rect 9938 908 10022 932
rect 9938 852 9952 908
rect 10008 852 10022 908
rect 9938 828 10022 852
rect 9938 772 9952 828
rect 10008 772 10022 828
rect 9938 748 10022 772
rect 9938 692 9952 748
rect 10008 692 10022 748
rect 9938 668 10022 692
rect 9938 612 9952 668
rect 10008 612 10022 668
rect 9938 588 10022 612
rect 9938 532 9952 588
rect 10008 532 10022 588
rect 9938 508 10022 532
rect 9938 452 9952 508
rect 10008 452 10022 508
rect 9938 428 10022 452
rect 9938 372 9952 428
rect 10008 372 10022 428
rect 9938 348 10022 372
rect 9938 292 9952 348
rect 10008 292 10022 348
rect 9938 268 10022 292
rect 9938 212 9952 268
rect 10008 212 10022 268
rect 9938 188 10022 212
rect 9938 132 9952 188
rect 10008 132 10022 188
rect 9938 108 10022 132
rect 9938 52 9952 108
rect 10008 52 10022 108
rect 9938 18 10022 52
<< via2 >>
rect 9952 4532 10008 4588
rect 9952 4452 10008 4508
rect 9952 4372 10008 4428
rect 9952 4292 10008 4348
rect 9952 4212 10008 4268
rect 9952 4132 10008 4188
rect 9952 4052 10008 4108
rect 9952 3972 10008 4028
rect 9952 3892 10008 3948
rect 9952 3812 10008 3868
rect 9952 3732 10008 3788
rect 9952 3652 10008 3708
rect 9952 3572 10008 3628
rect 9952 3492 10008 3548
rect 9952 3412 10008 3468
rect 9952 3332 10008 3388
rect 9952 3252 10008 3308
rect 9952 3172 10008 3228
rect 9952 3092 10008 3148
rect 9952 3012 10008 3068
rect 9952 2932 10008 2988
rect 9952 2852 10008 2908
rect 9952 2772 10008 2828
rect 9952 2692 10008 2748
rect 9952 2612 10008 2668
rect 9952 2532 10008 2588
rect 9952 2452 10008 2508
rect 9952 2372 10008 2428
rect 9952 2292 10008 2348
rect 9952 2212 10008 2268
rect 9952 2132 10008 2188
rect 9952 2052 10008 2108
rect 9952 1972 10008 2028
rect 9952 1892 10008 1948
rect 9952 1812 10008 1868
rect 9952 1732 10008 1788
rect 9952 1652 10008 1708
rect 9952 1572 10008 1628
rect 9952 1492 10008 1548
rect 9952 1412 10008 1468
rect 9952 1332 10008 1388
rect 9952 1252 10008 1308
rect 9952 1172 10008 1228
rect 9952 1092 10008 1148
rect 9952 1012 10008 1068
rect 9952 932 10008 988
rect 9952 852 10008 908
rect 9952 772 10008 828
rect 9952 692 10008 748
rect 9952 612 10008 668
rect 9952 532 10008 588
rect 9952 452 10008 508
rect 9952 372 10008 428
rect 9952 292 10008 348
rect 9952 212 10008 268
rect 9952 132 10008 188
rect 9952 52 10008 108
<< metal3 >>
rect 6000 5154 6320 5190
rect 6000 4930 6048 5154
rect 6272 4930 6320 5154
rect 6000 4640 6320 4930
rect 5016 4588 10032 4640
rect 5016 4532 9952 4588
rect 10008 4532 10032 4588
rect 5016 4508 10032 4532
rect 5016 4452 9952 4508
rect 10008 4452 10032 4508
rect 5016 4428 10032 4452
rect 5016 4374 9952 4428
rect 6000 4372 9952 4374
rect 10008 4372 10032 4428
rect 6000 4348 10032 4372
rect 6000 4292 9952 4348
rect 10008 4292 10032 4348
rect 6000 4268 10032 4292
rect 6000 4212 9952 4268
rect 10008 4212 10032 4268
rect 6000 4188 10032 4212
rect 6000 4132 9952 4188
rect 10008 4132 10032 4188
rect 6000 4108 10032 4132
rect 6000 4052 9952 4108
rect 10008 4052 10032 4108
rect 6000 4028 10032 4052
rect 6000 3972 9952 4028
rect 10008 3972 10032 4028
rect 6000 3948 10032 3972
rect 6000 3892 9952 3948
rect 10008 3892 10032 3948
rect 6000 3868 10032 3892
rect 6000 3812 9952 3868
rect 10008 3812 10032 3868
rect 6000 3788 10032 3812
rect 6000 3732 9952 3788
rect 10008 3732 10032 3788
rect 6000 3708 10032 3732
rect 6000 3652 9952 3708
rect 10008 3652 10032 3708
rect 6000 3628 10032 3652
rect 6000 3572 9952 3628
rect 10008 3572 10032 3628
rect 6000 3548 10032 3572
rect 6000 3492 9952 3548
rect 10008 3492 10032 3548
rect 6000 3468 10032 3492
rect 6000 3412 9952 3468
rect 10008 3412 10032 3468
rect 6000 3388 10032 3412
rect 6000 3332 9952 3388
rect 10008 3332 10032 3388
rect 6000 3308 10032 3332
rect 6000 3252 9952 3308
rect 10008 3252 10032 3308
rect 6000 3228 10032 3252
rect 6000 3172 9952 3228
rect 10008 3172 10032 3228
rect 6000 3148 10032 3172
rect 6000 3092 9952 3148
rect 10008 3092 10032 3148
rect 6000 3068 10032 3092
rect 6000 3012 9952 3068
rect 10008 3012 10032 3068
rect 6000 2988 10032 3012
rect 6000 2932 9952 2988
rect 10008 2932 10032 2988
rect 6000 2908 10032 2932
rect 6000 2852 9952 2908
rect 10008 2852 10032 2908
rect 6000 2828 10032 2852
rect 6000 2772 9952 2828
rect 10008 2772 10032 2828
rect 6000 2748 10032 2772
rect 6000 2692 9952 2748
rect 10008 2692 10032 2748
rect 6000 2668 10032 2692
rect 6000 2612 9952 2668
rect 10008 2612 10032 2668
rect 6000 2588 10032 2612
rect 6000 2532 9952 2588
rect 10008 2532 10032 2588
rect 6000 2508 10032 2532
rect 6000 2452 9952 2508
rect 10008 2452 10032 2508
rect 6000 2428 10032 2452
rect 6000 2372 9952 2428
rect 10008 2372 10032 2428
rect 6000 2348 10032 2372
rect 6000 2292 9952 2348
rect 10008 2292 10032 2348
rect 6000 2268 10032 2292
rect 6000 2212 9952 2268
rect 10008 2212 10032 2268
rect 6000 2188 10032 2212
rect 6000 2132 9952 2188
rect 10008 2132 10032 2188
rect 6000 2108 10032 2132
rect 6000 2052 9952 2108
rect 10008 2052 10032 2108
rect 6000 2028 10032 2052
rect 6000 1972 9952 2028
rect 10008 1972 10032 2028
rect 6000 1948 10032 1972
rect 6000 1892 9952 1948
rect 10008 1892 10032 1948
rect 6000 1868 10032 1892
rect 6000 1812 9952 1868
rect 10008 1812 10032 1868
rect 6000 1788 10032 1812
rect 6000 1732 9952 1788
rect 10008 1732 10032 1788
rect 6000 1708 10032 1732
rect 6000 1652 9952 1708
rect 10008 1652 10032 1708
rect 6000 1628 10032 1652
rect 6000 1572 9952 1628
rect 10008 1572 10032 1628
rect 6000 1548 10032 1572
rect 6000 1492 9952 1548
rect 10008 1492 10032 1548
rect 6000 1468 10032 1492
rect 6000 1412 9952 1468
rect 10008 1412 10032 1468
rect 6000 1388 10032 1412
rect 6000 1332 9952 1388
rect 10008 1332 10032 1388
rect 6000 1308 10032 1332
rect 6000 1252 9952 1308
rect 10008 1252 10032 1308
rect 6000 1228 10032 1252
rect 6000 1172 9952 1228
rect 10008 1172 10032 1228
rect 6000 1148 10032 1172
rect 6000 1092 9952 1148
rect 10008 1092 10032 1148
rect 6000 1068 10032 1092
rect 6000 1012 9952 1068
rect 10008 1012 10032 1068
rect 6000 988 10032 1012
rect 6000 932 9952 988
rect 10008 932 10032 988
rect 6000 908 10032 932
rect 6000 852 9952 908
rect 10008 852 10032 908
rect 6000 828 10032 852
rect 6000 772 9952 828
rect 10008 772 10032 828
rect 6000 748 10032 772
rect 6000 692 9952 748
rect 10008 692 10032 748
rect 6000 668 10032 692
rect 6000 612 9952 668
rect 10008 612 10032 668
rect 6000 588 10032 612
rect 6000 532 9952 588
rect 10008 532 10032 588
rect 6000 508 10032 532
rect 6000 452 9952 508
rect 10008 452 10032 508
rect 6000 428 10032 452
rect 6000 372 9952 428
rect 10008 372 10032 428
rect 6000 348 10032 372
rect 6000 292 9952 348
rect 10008 292 10032 348
rect 6000 268 10032 292
rect 6000 212 9952 268
rect 10008 212 10032 268
rect 6000 188 10032 212
rect 6000 132 9952 188
rect 10008 132 10032 188
rect 6000 108 10032 132
rect 6000 52 9952 108
rect 10008 52 10032 108
rect 4130 -116 4414 2
rect 6000 0 10032 52
rect 4130 -340 4162 -116
rect 4386 -340 4414 -116
rect 4130 -432 4414 -340
<< via3 >>
rect 6048 4930 6272 5154
rect 4162 -340 4386 -116
<< mimcap >>
rect 6100 4472 9860 4540
rect 6100 168 9656 4472
rect 9800 168 9860 4472
rect 6100 100 9860 168
<< mimcapcontact >>
rect 9656 168 9800 4472
<< metal4 >>
rect 8628 5268 9822 5306
rect 6000 5154 6320 5190
rect 3470 5094 4558 5142
rect 3470 4858 3506 5094
rect 3742 4858 4558 5094
rect 3470 4826 4558 4858
rect 4490 4498 4558 4826
rect 6000 4930 6048 5154
rect 6272 4930 6320 5154
rect 8848 5014 9822 5268
rect 6000 4640 6320 4930
rect 9634 4472 9822 5014
rect 9634 168 9656 4472
rect 9800 168 9822 4472
rect 9634 138 9822 168
rect 4130 -116 4414 2
rect 4130 -340 4162 -116
rect 4386 -340 4414 -116
rect 4130 -432 4414 -340
<< via4 >>
rect 3506 4858 3742 5094
rect 8612 5032 8848 5268
<< metal5 >>
rect 8526 5268 8936 5306
rect 3472 5094 3792 5140
rect 3472 4858 3506 5094
rect 3742 4858 3792 5094
rect 3472 4524 3792 4858
rect 8526 5032 8612 5268
rect 8848 5032 8936 5268
rect 3472 4500 3506 4524
rect 8526 4500 8936 5032
use sky130_fd_pr__cap_mim_m3_2_4SGG6N  sky130_fd_pr__cap_mim_m3_2_4SGG6N_0
timestamp 1640991954
transform 1 0 7323 0 1 2320
box -2231 -2321 2253 2321
use sky130_fd_pr__cap_mim_m3_1_9K4XRG  sky130_fd_pr__cap_mim_m3_1_9K4XRG_0
timestamp 1640991954
transform 1 0 4560 0 1 2320
box -456 -2320 456 2320
use sky130_fd_pr__cap_mim_m3_2_7PBNAZ  sky130_fd_pr__cap_mim_m3_2_7PBNAZ_0
timestamp 1640991954
transform 1 0 3739 0 1 2320
box -671 -2321 693 2321
<< labels >>
flabel metal4 s 6140 4764 6140 4764 0 FreeSans 2000 0 0 0 BOT
port 1 nsew
flabel metal4 s 4110 4986 4110 4986 0 FreeSans 2000 0 0 0 TOP_V
port 2 nsew
flabel metal4 s 9210 5152 9210 5152 0 FreeSans 2000 0 0 0 TOP_B
port 3 nsew
<< end >>
