magic
tech sky130A
magscale 1 2
timestamp 1641609411
<< nwell >>
rect 1366 442 2276 1080
<< pwell >>
rect 1376 -168 1882 432
<< nmos >>
rect 1566 32 1596 232
rect 1662 32 1692 232
<< pmos >>
rect 1566 662 1596 862
rect 1662 662 1692 862
rect 1758 662 1788 862
rect 1854 662 1884 862
rect 1950 662 1980 862
rect 2046 662 2076 862
<< ndiff >>
rect 1504 217 1566 232
rect 1504 183 1516 217
rect 1550 183 1566 217
rect 1504 149 1566 183
rect 1504 115 1516 149
rect 1550 115 1566 149
rect 1504 81 1566 115
rect 1504 47 1516 81
rect 1550 47 1566 81
rect 1504 32 1566 47
rect 1596 217 1662 232
rect 1596 183 1612 217
rect 1646 183 1662 217
rect 1596 149 1662 183
rect 1596 115 1612 149
rect 1646 115 1662 149
rect 1596 81 1662 115
rect 1596 47 1612 81
rect 1646 47 1662 81
rect 1596 32 1662 47
rect 1692 217 1754 232
rect 1692 183 1708 217
rect 1742 183 1754 217
rect 1692 149 1754 183
rect 1692 115 1708 149
rect 1742 115 1754 149
rect 1692 81 1754 115
rect 1692 47 1708 81
rect 1742 47 1754 81
rect 1692 32 1754 47
<< pdiff >>
rect 1504 845 1566 862
rect 1504 811 1516 845
rect 1550 811 1566 845
rect 1504 777 1566 811
rect 1504 743 1516 777
rect 1550 743 1566 777
rect 1504 709 1566 743
rect 1504 675 1516 709
rect 1550 675 1566 709
rect 1504 662 1566 675
rect 1596 845 1662 862
rect 1596 811 1612 845
rect 1646 811 1662 845
rect 1596 777 1662 811
rect 1596 743 1612 777
rect 1646 743 1662 777
rect 1596 709 1662 743
rect 1596 675 1612 709
rect 1646 675 1662 709
rect 1596 662 1662 675
rect 1692 845 1758 862
rect 1692 811 1708 845
rect 1742 811 1758 845
rect 1692 777 1758 811
rect 1692 743 1708 777
rect 1742 743 1758 777
rect 1692 709 1758 743
rect 1692 675 1708 709
rect 1742 675 1758 709
rect 1692 662 1758 675
rect 1788 845 1854 862
rect 1788 811 1804 845
rect 1838 811 1854 845
rect 1788 777 1854 811
rect 1788 743 1804 777
rect 1838 743 1854 777
rect 1788 709 1854 743
rect 1788 675 1804 709
rect 1838 675 1854 709
rect 1788 662 1854 675
rect 1884 845 1950 862
rect 1884 811 1900 845
rect 1934 811 1950 845
rect 1884 777 1950 811
rect 1884 743 1900 777
rect 1934 743 1950 777
rect 1884 709 1950 743
rect 1884 675 1900 709
rect 1934 675 1950 709
rect 1884 662 1950 675
rect 1980 845 2046 862
rect 1980 811 1996 845
rect 2030 811 2046 845
rect 1980 777 2046 811
rect 1980 743 1996 777
rect 2030 743 2046 777
rect 1980 709 2046 743
rect 1980 675 1996 709
rect 2030 675 2046 709
rect 1980 662 2046 675
rect 2076 845 2138 862
rect 2076 811 2092 845
rect 2126 811 2138 845
rect 2076 777 2138 811
rect 2076 743 2092 777
rect 2126 743 2138 777
rect 2076 709 2138 743
rect 2076 675 2092 709
rect 2126 675 2138 709
rect 2076 662 2138 675
<< ndiffc >>
rect 1516 183 1550 217
rect 1516 115 1550 149
rect 1516 47 1550 81
rect 1612 183 1646 217
rect 1612 115 1646 149
rect 1612 47 1646 81
rect 1708 183 1742 217
rect 1708 115 1742 149
rect 1708 47 1742 81
<< pdiffc >>
rect 1516 811 1550 845
rect 1516 743 1550 777
rect 1516 675 1550 709
rect 1612 811 1646 845
rect 1612 743 1646 777
rect 1612 675 1646 709
rect 1708 811 1742 845
rect 1708 743 1742 777
rect 1708 675 1742 709
rect 1804 811 1838 845
rect 1804 743 1838 777
rect 1804 675 1838 709
rect 1900 811 1934 845
rect 1900 743 1934 777
rect 1900 675 1934 709
rect 1996 811 2030 845
rect 1996 743 2030 777
rect 1996 675 2030 709
rect 2092 811 2126 845
rect 2092 743 2126 777
rect 2092 675 2126 709
<< psubdiff >>
rect 1402 372 1510 406
rect 1544 372 1578 406
rect 1612 372 1646 406
rect 1680 372 1714 406
rect 1748 372 1856 406
rect 1402 285 1436 372
rect 1402 217 1436 251
rect 1822 285 1856 372
rect 1402 149 1436 183
rect 1402 81 1436 115
rect 1402 13 1436 47
rect 1822 217 1856 251
rect 1822 149 1856 183
rect 1822 81 1856 115
rect 1822 13 1856 47
rect 1402 -108 1436 -21
rect 1822 -108 1856 -21
rect 1402 -142 1510 -108
rect 1544 -142 1578 -108
rect 1612 -142 1646 -108
rect 1680 -142 1714 -108
rect 1748 -142 1856 -108
<< nsubdiff >>
rect 1402 1010 1498 1044
rect 1532 1010 1566 1044
rect 1600 1010 1634 1044
rect 1668 1010 1702 1044
rect 1736 1010 1770 1044
rect 1804 1010 1838 1044
rect 1872 1010 1906 1044
rect 1940 1010 1974 1044
rect 2008 1010 2042 1044
rect 2076 1010 2110 1044
rect 2144 1010 2240 1044
rect 1402 948 1436 1010
rect 2206 948 2240 1010
rect 1402 880 1436 914
rect 2206 880 2240 914
rect 1402 812 1436 846
rect 1402 744 1436 778
rect 1402 676 1436 710
rect 2206 812 2240 846
rect 2206 744 2240 778
rect 2206 676 2240 710
rect 1402 608 1436 642
rect 1402 512 1436 574
rect 2206 608 2240 642
rect 2206 512 2240 574
rect 1402 478 1498 512
rect 1532 478 1566 512
rect 1600 478 1634 512
rect 1668 478 1702 512
rect 1736 478 1770 512
rect 1804 478 1838 512
rect 1872 478 1906 512
rect 1940 478 1974 512
rect 2008 478 2042 512
rect 2076 478 2110 512
rect 2144 478 2240 512
<< psubdiffcont >>
rect 1510 372 1544 406
rect 1578 372 1612 406
rect 1646 372 1680 406
rect 1714 372 1748 406
rect 1402 251 1436 285
rect 1822 251 1856 285
rect 1402 183 1436 217
rect 1402 115 1436 149
rect 1402 47 1436 81
rect 1822 183 1856 217
rect 1822 115 1856 149
rect 1822 47 1856 81
rect 1402 -21 1436 13
rect 1822 -21 1856 13
rect 1510 -142 1544 -108
rect 1578 -142 1612 -108
rect 1646 -142 1680 -108
rect 1714 -142 1748 -108
<< nsubdiffcont >>
rect 1498 1010 1532 1044
rect 1566 1010 1600 1044
rect 1634 1010 1668 1044
rect 1702 1010 1736 1044
rect 1770 1010 1804 1044
rect 1838 1010 1872 1044
rect 1906 1010 1940 1044
rect 1974 1010 2008 1044
rect 2042 1010 2076 1044
rect 2110 1010 2144 1044
rect 1402 914 1436 948
rect 1402 846 1436 880
rect 2206 914 2240 948
rect 1402 778 1436 812
rect 1402 710 1436 744
rect 1402 642 1436 676
rect 2206 846 2240 880
rect 2206 778 2240 812
rect 2206 710 2240 744
rect 1402 574 1436 608
rect 2206 642 2240 676
rect 2206 574 2240 608
rect 1498 478 1532 512
rect 1566 478 1600 512
rect 1634 478 1668 512
rect 1702 478 1736 512
rect 1770 478 1804 512
rect 1838 478 1872 512
rect 1906 478 1940 512
rect 1974 478 2008 512
rect 2042 478 2076 512
rect 2110 478 2144 512
<< poly >>
rect 1566 886 2076 916
rect 1566 862 1596 886
rect 1662 862 1692 886
rect 1758 862 1788 886
rect 1854 862 1884 886
rect 1950 862 1980 886
rect 2046 862 2076 886
rect 1566 636 1596 662
rect 1662 636 1692 662
rect 1758 636 1788 662
rect 1854 636 1884 662
rect 1950 636 1980 662
rect 2046 636 2076 662
rect 1566 630 2076 636
rect 1548 614 2076 630
rect 1548 580 1564 614
rect 1598 606 1756 614
rect 1598 580 1614 606
rect 1548 564 1614 580
rect 1740 580 1756 606
rect 1790 606 1948 614
rect 1790 580 1806 606
rect 1740 564 1806 580
rect 1932 580 1948 606
rect 1982 606 2076 614
rect 1982 580 1998 606
rect 1932 564 1998 580
rect 1644 304 1710 320
rect 1644 284 1660 304
rect 1566 270 1660 284
rect 1694 270 1710 304
rect 1566 254 1710 270
rect 1566 232 1596 254
rect 1662 232 1692 254
rect 1566 10 1596 32
rect 1662 10 1692 32
rect 1566 -20 1692 10
<< polycont >>
rect 1564 580 1598 614
rect 1756 580 1790 614
rect 1948 580 1982 614
rect 1660 270 1694 304
<< locali >>
rect 1402 1010 1498 1044
rect 1532 1010 1566 1044
rect 1600 1010 1634 1044
rect 1668 1010 1702 1044
rect 1736 1010 1770 1044
rect 1804 1010 1838 1044
rect 1872 1010 1906 1044
rect 1940 1010 1974 1044
rect 2008 1010 2042 1044
rect 2076 1010 2110 1044
rect 2144 1010 2240 1044
rect 1402 948 1436 1010
rect 1492 960 1550 976
rect 1526 926 1550 960
rect 1402 880 1436 914
rect 1402 812 1436 846
rect 1402 744 1436 778
rect 1402 676 1436 710
rect 1516 845 1550 926
rect 1516 777 1550 779
rect 1516 741 1550 743
rect 1516 656 1550 675
rect 1612 960 1646 976
rect 1646 926 2030 950
rect 1612 916 2030 926
rect 1612 845 1646 916
rect 1612 777 1646 811
rect 1612 709 1646 743
rect 1612 656 1646 675
rect 1708 845 1742 864
rect 1708 777 1742 779
rect 1708 741 1742 743
rect 1708 656 1742 675
rect 1804 845 1838 916
rect 1804 777 1838 811
rect 1804 709 1838 743
rect 1804 656 1838 675
rect 1900 845 1934 864
rect 1900 777 1934 779
rect 1900 741 1934 743
rect 1900 656 1934 675
rect 1996 845 2030 916
rect 2206 948 2240 1010
rect 2206 880 2240 914
rect 1996 777 2030 811
rect 1996 709 2030 743
rect 1996 656 2030 675
rect 2092 845 2126 864
rect 2092 777 2126 779
rect 2092 741 2126 743
rect 2092 656 2126 675
rect 2206 812 2240 846
rect 2206 744 2240 778
rect 2206 676 2240 710
rect 1402 608 1436 642
rect 2240 642 2326 672
rect 1548 580 1564 614
rect 1598 580 1614 614
rect 1740 580 1756 614
rect 1790 580 1806 614
rect 1932 580 1948 614
rect 1982 580 1998 614
rect 2206 608 2326 642
rect 1402 512 1436 574
rect 2240 574 2326 608
rect 2206 512 2326 574
rect 1402 478 1498 512
rect 1532 478 1566 512
rect 1600 478 1634 512
rect 1668 478 1702 512
rect 1736 478 1770 512
rect 1804 478 1838 512
rect 1872 478 1906 512
rect 1940 478 1974 512
rect 2008 478 2042 512
rect 2076 478 2110 512
rect 2144 492 2326 512
rect 2144 478 2240 492
rect 1402 372 1510 406
rect 1544 372 1578 406
rect 1612 372 1646 406
rect 1680 372 1714 406
rect 1748 372 1856 406
rect 1402 285 1436 372
rect 1822 362 1856 372
rect 1644 270 1660 304
rect 1694 270 1710 304
rect 1822 285 2326 362
rect 1402 217 1436 251
rect 1856 251 2326 285
rect 1402 149 1436 183
rect 1402 81 1436 115
rect 1402 13 1436 47
rect 1402 -108 1436 -21
rect 1516 217 1550 236
rect 1516 149 1550 151
rect 1516 113 1550 115
rect 1516 -22 1550 47
rect 1492 -38 1550 -22
rect 1526 -72 1550 -38
rect 1612 217 1646 236
rect 1612 149 1646 183
rect 1612 81 1646 115
rect 1612 -38 1646 47
rect 1708 217 1742 236
rect 1708 149 1742 151
rect 1708 113 1742 115
rect 1708 28 1742 47
rect 1822 217 2326 251
rect 1856 183 2326 217
rect 1822 182 2326 183
rect 1822 149 1856 182
rect 2706 134 2760 142
rect 1822 81 1856 115
rect 2706 100 2714 134
rect 2748 100 2760 134
rect 2706 92 2760 100
rect 1822 13 1856 47
rect 1822 -108 1856 -21
rect 1402 -142 1510 -108
rect 1544 -142 1578 -108
rect 1612 -142 1646 -108
rect 1680 -142 1714 -108
rect 1748 -142 1856 -108
<< viali >>
rect 1492 926 1526 960
rect 1516 811 1550 813
rect 1516 779 1550 811
rect 1516 709 1550 741
rect 1516 707 1550 709
rect 1612 926 1646 960
rect 1708 811 1742 813
rect 1708 779 1742 811
rect 1708 709 1742 741
rect 1708 707 1742 709
rect 1900 811 1934 813
rect 1900 779 1934 811
rect 1900 709 1934 741
rect 1900 707 1934 709
rect 2092 811 2126 813
rect 2092 779 2126 811
rect 2092 709 2126 741
rect 2092 707 2126 709
rect 1564 580 1598 614
rect 1756 580 1790 614
rect 1948 580 1982 614
rect 1660 270 1694 304
rect 1516 183 1550 185
rect 1516 151 1550 183
rect 1516 81 1550 113
rect 1516 79 1550 81
rect 1492 -72 1526 -38
rect 1708 183 1742 185
rect 1708 151 1742 183
rect 1708 81 1742 113
rect 1708 79 1742 81
rect 2284 100 2318 134
rect 2714 100 2748 134
rect 1612 -72 1646 -38
<< metal1 >>
rect 1476 969 1542 976
rect 1476 917 1483 969
rect 1535 917 1542 969
rect 1476 910 1542 917
rect 1596 969 1662 976
rect 1596 917 1603 969
rect 1655 917 1662 969
rect 1596 910 1662 917
rect 1516 860 2126 876
rect 1510 848 2132 860
rect 1510 813 1556 848
rect 1510 779 1516 813
rect 1550 779 1556 813
rect 1510 741 1556 779
rect 1510 707 1516 741
rect 1550 707 1556 741
rect 1510 660 1556 707
rect 1702 813 1748 848
rect 1702 779 1708 813
rect 1742 779 1748 813
rect 1702 741 1748 779
rect 1702 707 1708 741
rect 1742 707 1748 741
rect 1702 660 1748 707
rect 1894 813 1940 848
rect 1894 779 1900 813
rect 1934 779 1940 813
rect 1894 741 1940 779
rect 1894 707 1900 741
rect 1934 707 1940 741
rect 1894 660 1940 707
rect 2086 813 2132 848
rect 2086 779 2092 813
rect 2126 779 2132 813
rect 2086 741 2132 779
rect 2086 707 2092 741
rect 2126 707 2132 741
rect 2086 660 2132 707
rect 1552 614 2052 620
rect 1552 580 1564 614
rect 1598 580 1756 614
rect 1790 580 1948 614
rect 1982 580 2052 614
rect 1552 574 2052 580
rect 1994 452 2052 574
rect 1994 394 2882 452
rect 1644 304 2110 320
rect 1644 270 1660 304
rect 1694 270 2110 304
rect 1644 262 2110 270
rect 1510 185 1556 232
rect 1510 151 1516 185
rect 1550 151 1556 185
rect 1510 113 1556 151
rect 1510 79 1516 113
rect 1550 79 1556 113
rect 1510 44 1556 79
rect 1702 185 1748 232
rect 1702 151 1708 185
rect 1742 151 1748 185
rect 1702 113 1748 151
rect 1702 79 1708 113
rect 1742 79 1748 113
rect 2052 146 2110 262
rect 2824 146 2882 394
rect 2052 134 2330 146
rect 2052 100 2284 134
rect 2318 100 2330 134
rect 2052 88 2330 100
rect 2702 134 2882 146
rect 2702 100 2714 134
rect 2748 100 2882 134
rect 2702 86 2882 100
rect 1702 44 1748 79
rect 1510 32 1792 44
rect 1516 14 1792 32
rect 1476 -29 1542 -22
rect 1476 -81 1483 -29
rect 1535 -81 1542 -29
rect 1476 -88 1542 -81
rect 1596 -29 1662 -22
rect 1596 -81 1603 -29
rect 1655 -81 1662 -29
rect 1596 -88 1662 -81
<< via1 >>
rect 1483 960 1535 969
rect 1483 926 1492 960
rect 1492 926 1526 960
rect 1526 926 1535 960
rect 1483 917 1535 926
rect 1603 960 1655 969
rect 1603 926 1612 960
rect 1612 926 1646 960
rect 1646 926 1655 960
rect 1603 917 1655 926
rect 1483 -38 1535 -29
rect 1483 -72 1492 -38
rect 1492 -72 1526 -38
rect 1526 -72 1535 -38
rect 1483 -81 1535 -72
rect 1603 -38 1655 -29
rect 1603 -72 1612 -38
rect 1612 -72 1646 -38
rect 1646 -72 1655 -38
rect 1603 -81 1655 -72
<< metal2 >>
rect 1476 969 1544 976
rect 1476 917 1483 969
rect 1535 917 1544 969
rect 1476 -29 1544 917
rect 1476 -81 1483 -29
rect 1535 -81 1544 -29
rect 1476 -88 1544 -81
rect 1596 969 1662 976
rect 1596 917 1603 969
rect 1655 917 1662 969
rect 1596 -29 1662 917
rect 1596 -81 1603 -29
rect 1655 -81 1662 -29
rect 1596 -88 1662 -81
use INVMIN_v1p1  INVMIN_v1p1_0
timestamp 1641609411
transform 1 0 2576 0 1 192
box -300 -150 170 530
<< labels >>
flabel metal2 s 1508 940 1508 940 0 FreeSans 600 0 0 0 VIN
port 1 nsew
flabel metal2 s 1632 -54 1632 -54 0 FreeSans 600 0 0 0 VOUT
port 2 nsew
flabel metal1 s 1766 288 1766 288 0 FreeSans 600 0 0 0 CTR
port 3 nsew
flabel locali s 2296 588 2296 588 0 FreeSans 600 0 0 0 VDD
port 4 nsew
flabel locali s 2206 272 2206 272 0 FreeSans 600 0 0 0 VSS
port 5 nsew
<< end >>
