magic
tech sky130A
magscale 1 2
timestamp 1640975112
<< error_p >>
rect 14 -126 16 126
<< pwell >>
rect -98 -126 98 126
<< nmos >>
rect -14 -100 14 100
<< ndiff >>
rect -72 85 -14 100
rect -72 51 -60 85
rect -26 51 -14 85
rect -72 17 -14 51
rect -72 -17 -60 17
rect -26 -17 -14 17
rect -72 -51 -14 -17
rect -72 -85 -60 -51
rect -26 -85 -14 -51
rect -72 -100 -14 -85
rect 14 85 72 100
rect 14 51 26 85
rect 60 51 72 85
rect 14 17 72 51
rect 14 -17 26 17
rect 60 -17 72 17
rect 14 -51 72 -17
rect 14 -85 26 -51
rect 60 -85 72 -51
rect 14 -100 72 -85
<< ndiffc >>
rect -60 51 -26 85
rect -60 -17 -26 17
rect -60 -85 -26 -51
rect 26 51 60 85
rect 26 -17 60 17
rect 26 -85 60 -51
<< poly >>
rect -14 100 14 126
rect -14 -126 14 -100
<< locali >>
rect -60 85 -26 104
rect -60 17 -26 19
rect -60 -19 -26 -17
rect -60 -104 -26 -85
rect 26 85 60 104
rect 26 17 60 19
rect 26 -19 60 -17
rect 26 -104 60 -85
<< viali >>
rect -60 51 -26 53
rect -60 19 -26 51
rect -60 -51 -26 -19
rect -60 -53 -26 -51
rect 26 51 60 53
rect 26 19 60 51
rect 26 -51 60 -19
rect 26 -53 60 -51
<< metal1 >>
rect -66 53 -20 100
rect -66 19 -60 53
rect -26 19 -20 53
rect -66 -19 -20 19
rect -66 -53 -60 -19
rect -26 -53 -20 -19
rect -66 -100 -20 -53
rect 20 53 66 100
rect 20 19 26 53
rect 60 19 66 53
rect 20 -19 66 19
rect 20 -53 26 -19
rect 60 -53 66 -19
rect 20 -100 66 -53
<< end >>
