magic
tech sky130A
magscale 1 2
timestamp 1640975112
<< error_s >>
rect 22866 7800 23094 7827
rect 22894 7772 23094 7799
rect 22814 7701 22848 7765
rect 23079 7749 23094 7763
rect 23224 7749 23239 7763
rect 22864 7747 23094 7749
rect 23194 7748 23450 7749
rect 23224 7747 23450 7748
rect 23079 7703 23094 7719
rect 23224 7703 23239 7719
rect 22894 7667 23094 7694
rect 22894 7639 23094 7666
rect 22894 7600 23094 7627
rect 23224 7600 23451 7627
rect 22894 7572 23094 7599
rect 23225 7572 23423 7599
rect 22814 7501 22848 7565
rect 22864 7547 23120 7549
rect 23199 7547 23445 7549
rect 23098 7506 23132 7507
rect 23461 7501 23495 7565
rect 23225 7467 23423 7494
rect 23224 7439 23424 7466
rect 23224 7400 23424 7427
rect 23225 7372 23423 7399
rect 23199 7347 23445 7349
rect 23461 7301 23495 7365
rect 23225 7267 23423 7294
rect 20885 7246 21013 7247
rect 21077 7246 21205 7247
rect 21269 7246 21397 7247
rect 23224 7239 23424 7266
rect 23196 7227 23252 7228
rect 22856 7214 22928 7227
rect 22890 7194 22928 7214
rect 23196 7200 23424 7227
rect 23196 7199 23224 7200
rect 22814 7101 22848 7165
rect 22890 7160 22962 7193
rect 23196 7172 23424 7199
rect 22864 7148 23150 7149
rect 23168 7148 23450 7149
rect 22864 7147 23120 7148
rect 23198 7147 23450 7148
rect 22894 7067 23094 7094
rect 23224 7067 23424 7094
rect 22894 7039 23094 7066
rect 23224 7039 23424 7066
rect 22894 7000 23094 7027
rect 23224 7000 23424 7027
rect 22894 6972 23094 6999
rect 23224 6972 23424 6999
rect 22864 6948 23150 6949
rect 23168 6948 23450 6949
rect 22864 6947 23120 6948
rect 23198 6947 23450 6948
rect 22894 6867 22960 6894
rect 23196 6867 23424 6894
rect 23196 6866 23252 6867
rect 22894 6846 22932 6866
rect 22866 6839 22932 6846
rect 23224 6839 23424 6866
rect 23224 6838 23252 6839
rect 23224 6800 23424 6827
rect 23225 6772 23423 6799
rect 23199 6747 23445 6749
rect 23461 6701 23495 6765
rect 23225 6667 23423 6694
rect 23224 6639 23424 6666
rect 23224 6600 23424 6627
rect 23225 6572 23423 6599
rect 22814 6501 22848 6565
rect 22864 6547 23120 6549
rect 23199 6547 23445 6549
rect 23461 6501 23495 6565
rect 22894 6467 23094 6494
rect 23225 6467 23423 6494
rect 22894 6439 23094 6466
rect 23224 6439 23451 6466
rect 22894 6400 23094 6427
rect 22894 6372 23094 6399
rect 23079 6349 23094 6363
rect 23224 6349 23239 6363
rect 22864 6347 23094 6349
rect 23194 6348 23450 6349
rect 23224 6347 23450 6348
rect 23079 6303 23094 6319
rect 23224 6303 23239 6319
rect 22894 6267 23094 6294
rect 22866 6239 23094 6266
<< nwell >>
rect 20800 8076 20998 8234
rect 20734 7666 21644 8076
<< locali >>
rect 20866 7630 20884 7664
rect 20918 7630 20956 7664
rect 20990 7630 21028 7664
rect 21062 7630 21100 7664
rect 21134 7630 21172 7664
rect 21206 7630 21244 7664
rect 21278 7630 21316 7664
rect 21350 7630 21388 7664
rect 21422 7630 21460 7664
rect 21494 7630 21512 7664
rect 22756 7307 22816 7320
rect 22756 7273 22769 7307
rect 22803 7273 22816 7307
rect 22756 7260 22816 7273
rect 21874 6615 21934 6628
rect 21874 6581 21887 6615
rect 21921 6581 21934 6615
rect 21874 6568 21934 6581
rect 21224 6491 21284 6504
rect 21224 6457 21237 6491
rect 21271 6457 21284 6491
rect 21224 6444 21284 6457
<< viali >>
rect 20884 7630 20918 7664
rect 20956 7630 20990 7664
rect 21028 7630 21062 7664
rect 21100 7630 21134 7664
rect 21172 7630 21206 7664
rect 21244 7630 21278 7664
rect 21316 7630 21350 7664
rect 21388 7630 21422 7664
rect 21460 7630 21494 7664
rect 22769 7273 22803 7307
rect 21887 6581 21921 6615
rect 21237 6457 21271 6491
<< metal1 >>
rect 7826 9164 7920 9222
rect 22668 9130 23616 9242
rect 7778 7942 7862 7996
rect 20866 7676 21514 7848
rect 22122 7806 22774 8026
rect 20858 7664 21522 7676
rect 20858 7630 20884 7664
rect 20918 7630 20956 7664
rect 20990 7630 21028 7664
rect 21062 7630 21100 7664
rect 21134 7630 21172 7664
rect 21206 7630 21244 7664
rect 21278 7630 21316 7664
rect 21350 7630 21388 7664
rect 21422 7630 21460 7664
rect 21494 7630 21522 7664
rect 20858 7616 21522 7630
rect 23558 7564 23616 9130
rect 22744 7316 22828 7332
rect 22744 7264 22760 7316
rect 22812 7264 22828 7316
rect 22744 7248 22828 7264
rect 21862 6624 21946 6640
rect 21862 6572 21878 6624
rect 21930 6572 21946 6624
rect 21862 6556 21946 6572
rect 21212 6500 21298 6518
rect 21212 6448 21228 6500
rect 21280 6448 21298 6500
rect 21212 6430 21298 6448
rect 22122 6004 22774 6224
rect 23528 5874 23616 6444
rect 22106 5860 23616 5874
rect 22106 5808 22186 5860
rect 22238 5808 23616 5860
rect 22106 5794 23616 5808
<< via1 >>
rect 22760 7307 22812 7316
rect 22760 7273 22769 7307
rect 22769 7273 22803 7307
rect 22803 7273 22812 7307
rect 22760 7264 22812 7273
rect 21878 6615 21930 6624
rect 21878 6581 21887 6615
rect 21887 6581 21921 6615
rect 21921 6581 21930 6615
rect 21878 6572 21930 6581
rect 21228 6491 21280 6500
rect 21228 6457 21237 6491
rect 21237 6457 21271 6491
rect 21271 6457 21280 6491
rect 21228 6448 21280 6457
rect 22186 5808 22238 5860
<< metal2 >>
rect 9142 7660 9374 7780
rect 22022 7756 22246 8434
rect 22022 7692 22854 7756
rect 20790 7562 20912 7644
rect 20998 7513 21102 7562
rect 20998 7457 21021 7513
rect 21077 7457 21102 7513
rect 20998 7433 21102 7457
rect 20998 7377 21021 7433
rect 21077 7377 21102 7433
rect 20998 7353 21102 7377
rect 20998 7297 21021 7353
rect 21077 7297 21102 7353
rect 20998 7273 21102 7297
rect 20998 7217 21021 7273
rect 21077 7217 21102 7273
rect 20998 7193 21102 7217
rect 20998 7137 21021 7193
rect 21077 7137 21102 7193
rect 20998 7113 21102 7137
rect 20998 7057 21021 7113
rect 21077 7057 21102 7113
rect 20998 7046 21102 7057
rect 22402 7316 22822 7328
rect 22402 7264 22760 7316
rect 22812 7264 22822 7316
rect 22402 7254 22822 7264
rect 22402 6636 22476 7254
rect 21868 6624 22476 6636
rect 21868 6572 21878 6624
rect 21930 6572 22476 6624
rect 21868 6562 22476 6572
rect 21218 6500 22248 6510
rect 21218 6448 21228 6500
rect 21280 6448 22248 6500
rect 21218 6438 22248 6448
rect 22176 5860 22248 6438
rect 22176 5808 22186 5860
rect 22238 5808 22248 5860
rect 22176 5798 22248 5808
rect 22994 5626 23062 6528
rect 22220 5472 23062 5626
<< via2 >>
rect 21021 7457 21077 7513
rect 21021 7377 21077 7433
rect 21021 7297 21077 7353
rect 21021 7217 21077 7273
rect 21021 7137 21077 7193
rect 21021 7057 21077 7113
<< metal3 >>
rect 20998 7513 21102 7562
rect 20998 7477 21021 7513
rect 21077 7477 21102 7513
rect 20998 7413 21017 7477
rect 21081 7413 21102 7477
rect 20998 7397 21021 7413
rect 21077 7397 21102 7413
rect 20998 7333 21017 7397
rect 21081 7333 21102 7397
rect 20998 7317 21021 7333
rect 21077 7317 21102 7333
rect 20998 7253 21017 7317
rect 21081 7253 21102 7317
rect 20998 7237 21021 7253
rect 21077 7237 21102 7253
rect 20998 7173 21017 7237
rect 21081 7173 21102 7237
rect 20998 7157 21021 7173
rect 21077 7157 21102 7173
rect 20998 7093 21017 7157
rect 21081 7093 21102 7157
rect 20998 7057 21021 7093
rect 21077 7057 21102 7093
rect 20998 7046 21102 7057
<< via3 >>
rect 21017 7457 21021 7477
rect 21021 7457 21077 7477
rect 21077 7457 21081 7477
rect 21017 7433 21081 7457
rect 21017 7413 21021 7433
rect 21021 7413 21077 7433
rect 21077 7413 21081 7433
rect 21017 7377 21021 7397
rect 21021 7377 21077 7397
rect 21077 7377 21081 7397
rect 21017 7353 21081 7377
rect 21017 7333 21021 7353
rect 21021 7333 21077 7353
rect 21077 7333 21081 7353
rect 21017 7297 21021 7317
rect 21021 7297 21077 7317
rect 21077 7297 21081 7317
rect 21017 7273 21081 7297
rect 21017 7253 21021 7273
rect 21021 7253 21077 7273
rect 21077 7253 21081 7273
rect 21017 7217 21021 7237
rect 21021 7217 21077 7237
rect 21077 7217 21081 7237
rect 21017 7193 21081 7217
rect 21017 7173 21021 7193
rect 21021 7173 21077 7193
rect 21077 7173 21081 7193
rect 21017 7137 21021 7157
rect 21021 7137 21077 7157
rect 21077 7137 21081 7157
rect 21017 7113 21081 7137
rect 21017 7093 21021 7113
rect 21021 7093 21077 7113
rect 21077 7093 21081 7113
<< metal4 >>
rect 20620 8356 21102 8502
rect 20420 8320 21102 8356
rect 20998 7477 21102 8320
rect 20998 7413 21017 7477
rect 21081 7413 21102 7477
rect 20998 7397 21102 7413
rect 20998 7333 21017 7397
rect 21081 7333 21102 7397
rect 20998 7317 21102 7333
rect 20998 7253 21017 7317
rect 21081 7253 21102 7317
rect 20998 7237 21102 7253
rect 20998 7173 21017 7237
rect 21081 7173 21102 7237
rect 20998 7157 21102 7173
rect 20998 7093 21017 7157
rect 21081 7093 21102 7157
rect 20998 7046 21102 7093
<< via4 >>
rect 20384 8356 20620 8592
<< metal5 >>
rect 20280 8592 20514 8676
rect 20280 8356 20384 8592
rect 20620 8356 20654 8504
rect 20280 8320 20654 8356
rect 20654 5208 21574 5528
use OSC_v3p2  OSC_v3p2_1
timestamp 1640975112
transform 1 0 1718 0 -1 14404
box -12 10 20956 6760
use OSC_v3p2  OSC_v3p2_0
timestamp 1640975112
transform 1 0 1718 0 1 -374
box -12 10 20956 6760
use DFF_v3p1  DFF_v3p1_0
timestamp 1640975112
transform 0 -1 23450 1 0 6860
box -678 -204 986 904
use PASSGATE_v1p1  PASSGATE_v1p1_0
timestamp 1640975112
transform 1 0 19368 0 1 6586
box 1366 -168 2882 1080
<< labels >>
flabel metal1 s 7808 7968 7808 7968 0 FreeSans 2000 0 0 0 VDD
port 1 nsew
flabel metal1 s 7874 9190 7874 9190 0 FreeSans 2000 0 0 0 VSS
port 2 nsew
flabel metal2 s 9244 7732 9244 7732 0 FreeSans 2000 0 0 0 SENS_IN
port 3 nsew
flabel metal5 s 20956 5398 20956 5398 0 FreeSans 2000 0 0 0 REF_IN
port 4 nsew
flabel metal2 s 22458 7288 22458 7288 0 FreeSans 2000 0 0 0 DOUT
port 5 nsew
<< end >>
