magic
tech sky130A
magscale 1 2
timestamp 1640991954
<< locali >>
rect 19462 5928 19674 6028
rect 19462 5822 19515 5928
rect 19621 5822 19674 5928
rect 20304 5982 20528 6028
rect 20304 5876 20363 5982
rect 20469 5876 20528 5982
rect 20304 5846 20528 5876
rect 19462 5802 19674 5822
<< viali >>
rect 19515 5822 19621 5928
rect 20363 5876 20469 5982
<< metal1 >>
rect 19112 6486 19464 6558
rect 5000 6374 19464 6486
rect 19112 6372 19464 6374
rect 19464 6046 20404 6068
rect 19464 6044 20092 6046
rect 19462 5928 19674 5950
rect 19462 5901 19515 5928
rect 19621 5901 19674 5928
rect 19462 5849 19510 5901
rect 19626 5849 19674 5901
rect 19462 5822 19515 5849
rect 19621 5822 19674 5849
rect 19462 5802 19674 5822
rect 19776 5270 20092 6044
rect 20304 5982 20528 6000
rect 20304 5955 20363 5982
rect 20469 5955 20528 5982
rect 20304 5903 20358 5955
rect 20474 5903 20528 5955
rect 20304 5876 20363 5903
rect 20469 5876 20528 5903
rect 20304 5846 20528 5876
rect 19776 5268 20404 5270
rect 4722 5168 20956 5268
<< via1 >>
rect 19510 5849 19515 5901
rect 19515 5849 19562 5901
rect 19574 5849 19621 5901
rect 19621 5849 19626 5901
rect 20358 5903 20363 5955
rect 20363 5903 20410 5955
rect 20422 5903 20469 5955
rect 20469 5903 20474 5955
<< metal2 >>
rect 3964 6592 19294 6760
rect 3964 5508 4132 6592
rect 5126 5504 11132 5676
rect 12126 5504 18132 5676
rect 19126 5504 19294 6592
rect 20304 5955 20528 6000
rect 19462 5901 19674 5950
rect 19462 5849 19510 5901
rect 19562 5849 19574 5901
rect 19626 5849 19674 5901
rect 19462 5802 19674 5849
rect 20304 5903 20358 5955
rect 20410 5903 20422 5955
rect 20474 5903 20528 5955
rect 20304 5846 20528 5903
rect 17960 5362 18132 5504
rect 19502 5362 19674 5802
rect 17958 5190 19676 5362
<< metal3 >>
rect 2840 5002 3000 5162
rect 9840 5002 10000 5162
rect 16840 5002 17000 5162
<< metal5 >>
rect 392 5582 5856 5902
rect 7392 5582 12856 5902
rect 14392 5582 18936 5902
use INVandCAP_v1p1  INVandCAP_v1p1_0
timestamp 1640991954
transform 1 0 13988 0 1 10
box 0 0 6968 6476
use INVandCAP_v1p1  INVandCAP_v1p1_1
timestamp 1640991954
transform 1 0 6988 0 1 10
box 0 0 6968 6476
use INVandCAP_v1p1  INVandCAP_v1p1_2
timestamp 1640991954
transform 1 0 -12 0 1 10
box 0 0 6968 6476
use BUFFMIN_v1p1  BUFFMIN_v1p1_0
timestamp 1640991954
transform 1 0 19494 0 1 5938
box -30 -10 910 670
<< labels >>
flabel metal1 s 5626 6424 5626 6424 0 FreeSans 2000 0 0 0 VDD
port 1 nsew
flabel metal1 s 5512 5204 5512 5204 0 FreeSans 2000 0 0 0 VSS
port 2 nsew
flabel metal2 s 4048 6666 4048 6666 0 FreeSans 2000 0 0 0 SENS_IN
port 3 nsew
flabel metal2 s 7040 5580 7040 5580 0 FreeSans 2000 0 0 0 N1
port 4 nsew
flabel metal5 s 16012 5754 16012 5754 0 FreeSans 2000 0 0 0 CON_CV
port 5 nsew
flabel locali s 20362 6000 20362 6000 0 FreeSans 2000 0 0 0 N2
port 6 nsew
<< end >>
