magic
tech sky130A
magscale 1 2
timestamp 1640991954
<< metal4 >>
rect -2231 2198 2231 2320
rect -2231 1962 1975 2198
rect 2211 1962 2231 2198
rect -2231 1878 2231 1962
rect -2231 1642 1975 1878
rect 2211 1642 2231 1878
rect -2231 1558 2231 1642
rect -2231 1322 1975 1558
rect 2211 1322 2231 1558
rect -2231 1238 2231 1322
rect -2231 1002 1975 1238
rect 2211 1002 2231 1238
rect -2231 918 2231 1002
rect -2231 682 1975 918
rect 2211 682 2231 918
rect -2231 598 2231 682
rect -2231 362 1975 598
rect 2211 362 2231 598
rect -2231 278 2231 362
rect -2231 42 1975 278
rect 2211 42 2231 278
rect -2231 -42 2231 42
rect -2231 -278 1975 -42
rect 2211 -278 2231 -42
rect -2231 -362 2231 -278
rect -2231 -598 1975 -362
rect 2211 -598 2231 -362
rect -2231 -682 2231 -598
rect -2231 -918 1975 -682
rect 2211 -918 2231 -682
rect -2231 -1002 2231 -918
rect -2231 -1238 1975 -1002
rect 2211 -1238 2231 -1002
rect -2231 -1322 2231 -1238
rect -2231 -1558 1975 -1322
rect 2211 -1558 2231 -1322
rect -2231 -1642 2231 -1558
rect -2231 -1878 1975 -1642
rect 2211 -1878 2231 -1642
rect -2231 -1962 2231 -1878
rect -2231 -2198 1975 -1962
rect 2211 -2198 2231 -1962
rect -2231 -2320 2231 -2198
<< via4 >>
rect 1975 1962 2211 2198
rect 1975 1642 2211 1878
rect 1975 1322 2211 1558
rect 1975 1002 2211 1238
rect 1975 682 2211 918
rect 1975 362 2211 598
rect 1975 42 2211 278
rect 1975 -278 2211 -42
rect 1975 -598 2211 -362
rect 1975 -918 2211 -682
rect 1975 -1238 2211 -1002
rect 1975 -1558 2211 -1322
rect 1975 -1878 2211 -1642
rect 1975 -2198 2211 -1962
<< mimcap2 >>
rect -2131 2038 1629 2220
rect -2131 -2038 -1969 2038
rect 1467 -2038 1629 2038
rect -2131 -2220 1629 -2038
<< mimcap2contact >>
rect -1969 -2038 1467 2038
<< metal5 >>
rect -2115 2038 1613 2204
rect -2115 -2038 -1969 2038
rect 1467 -2038 1613 2038
rect -2115 -2204 1613 -2038
rect 1933 2198 2253 2321
rect 1933 1962 1975 2198
rect 2211 1962 2253 2198
rect 1933 1878 2253 1962
rect 1933 1642 1975 1878
rect 2211 1642 2253 1878
rect 1933 1558 2253 1642
rect 1933 1322 1975 1558
rect 2211 1322 2253 1558
rect 1933 1238 2253 1322
rect 1933 1002 1975 1238
rect 2211 1002 2253 1238
rect 1933 918 2253 1002
rect 1933 682 1975 918
rect 2211 682 2253 918
rect 1933 598 2253 682
rect 1933 362 1975 598
rect 2211 362 2253 598
rect 1933 278 2253 362
rect 1933 42 1975 278
rect 2211 42 2253 278
rect 1933 -42 2253 42
rect 1933 -278 1975 -42
rect 2211 -278 2253 -42
rect 1933 -362 2253 -278
rect 1933 -598 1975 -362
rect 2211 -598 2253 -362
rect 1933 -682 2253 -598
rect 1933 -918 1975 -682
rect 2211 -918 2253 -682
rect 1933 -1002 2253 -918
rect 1933 -1238 1975 -1002
rect 2211 -1238 2253 -1002
rect 1933 -1322 2253 -1238
rect 1933 -1558 1975 -1322
rect 2211 -1558 2253 -1322
rect 1933 -1642 2253 -1558
rect 1933 -1878 1975 -1642
rect 2211 -1878 2253 -1642
rect 1933 -1962 2253 -1878
rect 1933 -2198 1975 -1962
rect 2211 -2198 2253 -1962
rect 1933 -2321 2253 -2198
<< properties >>
string FIXED_BBOX -2231 -2320 1729 2320
<< end >>
