magic
tech sky130A
magscale 1 2
timestamp 1641609411
<< nwell >>
rect 20800 8076 20998 8234
rect 20734 7666 21644 8076
<< locali >>
rect 20866 7630 20884 7664
rect 20918 7630 20956 7664
rect 20990 7630 21028 7664
rect 21062 7630 21100 7664
rect 21134 7630 21172 7664
rect 21206 7630 21244 7664
rect 21278 7630 21316 7664
rect 21350 7630 21388 7664
rect 21422 7630 21460 7664
rect 21494 7630 21512 7664
rect 22756 7307 22816 7320
rect 22756 7273 22769 7307
rect 22803 7273 22816 7307
rect 22756 7244 22816 7273
rect 21874 6615 21934 6628
rect 21874 6581 21887 6615
rect 21921 6581 21934 6615
rect 21874 6568 21934 6581
rect 21224 6491 21284 6504
rect 21224 6457 21237 6491
rect 21271 6457 21284 6491
rect 21224 6444 21284 6457
<< viali >>
rect 20884 7630 20918 7664
rect 20956 7630 20990 7664
rect 21028 7630 21062 7664
rect 21100 7630 21134 7664
rect 21172 7630 21206 7664
rect 21244 7630 21278 7664
rect 21316 7630 21350 7664
rect 21388 7630 21422 7664
rect 21460 7630 21494 7664
rect 22769 7273 22803 7307
rect 21887 6581 21921 6615
rect 21237 6457 21271 6491
<< metal1 >>
rect 7826 9164 7920 9222
rect 22668 9130 23616 9242
rect 7778 7942 7862 7996
rect 20866 7676 21514 7848
rect 22122 7806 22774 8026
rect 23558 7818 23616 9130
rect 22788 7750 22864 7766
rect 22788 7698 22795 7750
rect 22847 7698 22864 7750
rect 22788 7692 22864 7698
rect 20858 7664 21522 7676
rect 20858 7630 20884 7664
rect 20918 7630 20956 7664
rect 20990 7630 21028 7664
rect 21062 7630 21100 7664
rect 21134 7630 21172 7664
rect 21206 7630 21244 7664
rect 21278 7630 21316 7664
rect 21350 7630 21388 7664
rect 21422 7630 21460 7664
rect 21494 7630 21522 7664
rect 20858 7616 21522 7630
rect 23558 7658 23638 7818
rect 23558 7600 23616 7658
rect 23558 7564 23638 7600
rect 22744 7316 22828 7332
rect 22744 7264 22760 7316
rect 22812 7264 22828 7316
rect 22744 7248 22828 7264
rect 21862 6624 21946 6640
rect 21862 6572 21878 6624
rect 21930 6572 21946 6624
rect 21862 6556 21946 6572
rect 21212 6500 21298 6518
rect 21212 6448 21228 6500
rect 21280 6448 21298 6500
rect 21212 6430 21298 6448
rect 23528 6408 23616 6444
rect 23528 6248 23638 6408
rect 22590 6224 23094 6232
rect 22122 6004 23094 6224
rect 23528 5874 23616 6248
rect 22106 5860 23616 5874
rect 22106 5808 22186 5860
rect 22238 5808 23616 5860
rect 22106 5794 23616 5808
<< via1 >>
rect 22795 7698 22847 7750
rect 22760 7307 22812 7316
rect 22760 7273 22769 7307
rect 22769 7273 22803 7307
rect 22803 7273 22812 7307
rect 22760 7264 22812 7273
rect 21878 6615 21930 6624
rect 21878 6581 21887 6615
rect 21887 6581 21921 6615
rect 21921 6581 21930 6615
rect 21878 6572 21930 6581
rect 21228 6491 21280 6500
rect 21228 6457 21237 6491
rect 21237 6457 21271 6491
rect 21271 6457 21280 6491
rect 21228 6448 21280 6457
rect 22186 5808 22238 5860
<< metal2 >>
rect 9142 7660 9374 7780
rect 22022 7756 22246 8434
rect 22022 7750 22854 7756
rect 22022 7698 22795 7750
rect 22847 7698 22854 7750
rect 22022 7692 22854 7698
rect 20790 7562 20912 7644
rect 20998 7513 21102 7562
rect 20998 7457 21021 7513
rect 21077 7457 21102 7513
rect 20998 7433 21102 7457
rect 20998 7377 21021 7433
rect 21077 7377 21102 7433
rect 20998 7353 21102 7377
rect 20998 7297 21021 7353
rect 21077 7297 21102 7353
rect 20998 7273 21102 7297
rect 20998 7217 21021 7273
rect 21077 7217 21102 7273
rect 20998 7193 21102 7217
rect 20998 7137 21021 7193
rect 21077 7137 21102 7193
rect 20998 7113 21102 7137
rect 20998 7057 21021 7113
rect 21077 7057 21102 7113
rect 20998 7046 21102 7057
rect 22402 7316 22822 7328
rect 22402 7264 22760 7316
rect 22812 7264 22822 7316
rect 22402 7254 22822 7264
rect 22402 6636 22476 7254
rect 21868 6624 22476 6636
rect 21868 6572 21878 6624
rect 21930 6572 22476 6624
rect 21868 6562 22476 6572
rect 21218 6500 22248 6510
rect 21218 6448 21228 6500
rect 21280 6448 22248 6500
rect 21218 6438 22248 6448
rect 22176 5860 22248 6438
rect 22176 5808 22186 5860
rect 22238 5808 22248 5860
rect 22176 5798 22248 5808
rect 22994 5626 23062 6528
rect 22220 5472 23062 5626
<< via2 >>
rect 21021 7457 21077 7513
rect 21021 7377 21077 7433
rect 21021 7297 21077 7353
rect 21021 7217 21077 7273
rect 21021 7137 21077 7193
rect 21021 7057 21077 7113
<< metal3 >>
rect 20998 7513 21102 7562
rect 20998 7477 21021 7513
rect 21077 7477 21102 7513
rect 20998 7413 21017 7477
rect 21081 7413 21102 7477
rect 20998 7397 21021 7413
rect 21077 7397 21102 7413
rect 20998 7333 21017 7397
rect 21081 7333 21102 7397
rect 20998 7317 21021 7333
rect 21077 7317 21102 7333
rect 20998 7253 21017 7317
rect 21081 7253 21102 7317
rect 20998 7237 21021 7253
rect 21077 7237 21102 7253
rect 20998 7173 21017 7237
rect 21081 7173 21102 7237
rect 20998 7157 21021 7173
rect 21077 7157 21102 7173
rect 20998 7093 21017 7157
rect 21081 7093 21102 7157
rect 20998 7057 21021 7093
rect 21077 7057 21102 7093
rect 20998 7046 21102 7057
<< via3 >>
rect 21017 7457 21021 7477
rect 21021 7457 21077 7477
rect 21077 7457 21081 7477
rect 21017 7433 21081 7457
rect 21017 7413 21021 7433
rect 21021 7413 21077 7433
rect 21077 7413 21081 7433
rect 21017 7377 21021 7397
rect 21021 7377 21077 7397
rect 21077 7377 21081 7397
rect 21017 7353 21081 7377
rect 21017 7333 21021 7353
rect 21021 7333 21077 7353
rect 21077 7333 21081 7353
rect 21017 7297 21021 7317
rect 21021 7297 21077 7317
rect 21077 7297 21081 7317
rect 21017 7273 21081 7297
rect 21017 7253 21021 7273
rect 21021 7253 21077 7273
rect 21077 7253 21081 7273
rect 21017 7217 21021 7237
rect 21021 7217 21077 7237
rect 21077 7217 21081 7237
rect 21017 7193 21081 7217
rect 21017 7173 21021 7193
rect 21021 7173 21077 7193
rect 21077 7173 21081 7193
rect 21017 7137 21021 7157
rect 21021 7137 21077 7157
rect 21077 7137 21081 7157
rect 21017 7113 21081 7137
rect 21017 7093 21021 7113
rect 21021 7093 21077 7113
rect 21077 7093 21081 7113
<< metal4 >>
rect 20620 8356 21102 8502
rect 20420 8320 21102 8356
rect 20998 7477 21102 8320
rect 20998 7413 21017 7477
rect 21081 7413 21102 7477
rect 20998 7397 21102 7413
rect 20998 7333 21017 7397
rect 21081 7333 21102 7397
rect 20998 7317 21102 7333
rect 20998 7253 21017 7317
rect 21081 7253 21102 7317
rect 20998 7237 21102 7253
rect 20998 7173 21017 7237
rect 21081 7173 21102 7237
rect 20998 7157 21102 7173
rect 20998 7093 21017 7157
rect 21081 7093 21102 7157
rect 20998 7046 21102 7093
<< via4 >>
rect 20384 8356 20620 8592
<< metal5 >>
rect 20280 8592 20514 8676
rect 20280 8356 20384 8592
rect 20620 8356 20654 8504
rect 20280 8320 20654 8356
rect 20654 5208 21574 5528
use PASSGATE_v1p2  PASSGATE_v1p2_0
timestamp 1641609411
transform 1 0 19368 0 1 6586
box 1366 -168 2882 1080
use DFF_v4p1  DFF_v4p1_0
timestamp 1641609411
transform 0 -1 23156 1 0 6824
box -636 -644 1036 626
use OSC_v3p2  OSC_v3p2_0 ~/Documents/Postdoc/github/caravel_user_project_analog/mag
timestamp 1641609411
transform 1 0 1718 0 -1 14404
box -12 10 20956 6760
use OSC_v3p2  OSC_v3p2_1
timestamp 1641609411
transform 1 0 1718 0 1 -374
box -12 10 20956 6760
<< labels >>
flabel metal1 s 7808 7968 7808 7968 0 FreeSans 2000 0 0 0 VDD
port 1 nsew
flabel metal1 s 7874 9190 7874 9190 0 FreeSans 2000 0 0 0 VSS
port 2 nsew
flabel metal2 s 9244 7732 9244 7732 0 FreeSans 2000 0 0 0 SENS_IN
port 3 nsew
flabel metal5 s 20956 5398 20956 5398 0 FreeSans 2000 0 0 0 REF_IN
port 4 nsew
flabel metal2 s 22458 7288 22458 7288 0 FreeSans 2000 0 0 0 DOUT
port 5 nsew
<< end >>
