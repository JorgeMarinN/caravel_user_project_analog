magic
tech sky130A
magscale 1 2
timestamp 1640975112
<< nwell >>
rect 1366 442 2276 1080
<< pwell >>
rect 1376 -168 1882 432
<< nmos >>
rect 1566 32 1596 232
rect 1662 32 1692 232
<< pmos >>
rect 1566 661 1596 861
rect 1662 661 1692 861
rect 1758 661 1788 861
rect 1854 661 1884 861
rect 1950 661 1980 861
rect 2046 661 2076 861
<< ndiff >>
rect 1504 217 1566 232
rect 1504 183 1516 217
rect 1550 183 1566 217
rect 1504 149 1566 183
rect 1504 115 1516 149
rect 1550 115 1566 149
rect 1504 81 1566 115
rect 1504 47 1516 81
rect 1550 47 1566 81
rect 1504 32 1566 47
rect 1596 217 1662 232
rect 1596 183 1612 217
rect 1646 183 1662 217
rect 1596 149 1662 183
rect 1596 115 1612 149
rect 1646 115 1662 149
rect 1596 81 1662 115
rect 1596 47 1612 81
rect 1646 47 1662 81
rect 1596 32 1662 47
rect 1692 217 1754 232
rect 1692 183 1708 217
rect 1742 183 1754 217
rect 1692 149 1754 183
rect 1692 115 1708 149
rect 1742 115 1754 149
rect 1692 81 1754 115
rect 1692 47 1708 81
rect 1742 47 1754 81
rect 1692 32 1754 47
<< pdiff >>
rect 1504 846 1566 861
rect 1504 812 1516 846
rect 1550 812 1566 846
rect 1504 778 1566 812
rect 1504 744 1516 778
rect 1550 744 1566 778
rect 1504 710 1566 744
rect 1504 676 1516 710
rect 1550 676 1566 710
rect 1504 661 1566 676
rect 1596 846 1662 861
rect 1596 812 1612 846
rect 1646 812 1662 846
rect 1596 778 1662 812
rect 1596 744 1612 778
rect 1646 744 1662 778
rect 1596 710 1662 744
rect 1596 676 1612 710
rect 1646 676 1662 710
rect 1596 661 1662 676
rect 1692 846 1758 861
rect 1692 812 1708 846
rect 1742 812 1758 846
rect 1692 778 1758 812
rect 1692 744 1708 778
rect 1742 744 1758 778
rect 1692 710 1758 744
rect 1692 676 1708 710
rect 1742 676 1758 710
rect 1692 661 1758 676
rect 1788 846 1854 861
rect 1788 812 1804 846
rect 1838 812 1854 846
rect 1788 778 1854 812
rect 1788 744 1804 778
rect 1838 744 1854 778
rect 1788 710 1854 744
rect 1788 676 1804 710
rect 1838 676 1854 710
rect 1788 661 1854 676
rect 1884 846 1950 861
rect 1884 812 1900 846
rect 1934 812 1950 846
rect 1884 778 1950 812
rect 1884 744 1900 778
rect 1934 744 1950 778
rect 1884 710 1950 744
rect 1884 676 1900 710
rect 1934 676 1950 710
rect 1884 661 1950 676
rect 1980 846 2046 861
rect 1980 812 1996 846
rect 2030 812 2046 846
rect 1980 778 2046 812
rect 1980 744 1996 778
rect 2030 744 2046 778
rect 1980 710 2046 744
rect 1980 676 1996 710
rect 2030 676 2046 710
rect 1980 661 2046 676
rect 2076 846 2138 861
rect 2076 812 2092 846
rect 2126 812 2138 846
rect 2076 778 2138 812
rect 2076 744 2092 778
rect 2126 744 2138 778
rect 2076 710 2138 744
rect 2076 676 2092 710
rect 2126 676 2138 710
rect 2076 661 2138 676
<< ndiffc >>
rect 1516 183 1550 217
rect 1516 115 1550 149
rect 1516 47 1550 81
rect 1612 183 1646 217
rect 1612 115 1646 149
rect 1612 47 1646 81
rect 1708 183 1742 217
rect 1708 115 1742 149
rect 1708 47 1742 81
<< pdiffc >>
rect 1516 812 1550 846
rect 1516 744 1550 778
rect 1516 676 1550 710
rect 1612 812 1646 846
rect 1612 744 1646 778
rect 1612 676 1646 710
rect 1708 812 1742 846
rect 1708 744 1742 778
rect 1708 676 1742 710
rect 1804 812 1838 846
rect 1804 744 1838 778
rect 1804 676 1838 710
rect 1900 812 1934 846
rect 1900 744 1934 778
rect 1900 676 1934 710
rect 1996 812 2030 846
rect 1996 744 2030 778
rect 1996 676 2030 710
rect 2092 812 2126 846
rect 2092 744 2126 778
rect 2092 676 2126 710
<< psubdiff >>
rect 1402 372 1510 406
rect 1544 372 1578 406
rect 1612 372 1646 406
rect 1680 372 1714 406
rect 1748 372 1856 406
rect 1402 285 1436 372
rect 1402 217 1436 251
rect 1822 285 1856 372
rect 1402 149 1436 183
rect 1402 81 1436 115
rect 1402 13 1436 47
rect 1822 217 1856 251
rect 1822 149 1856 183
rect 1822 81 1856 115
rect 1822 13 1856 47
rect 1402 -108 1436 -21
rect 1822 -108 1856 -21
rect 1402 -142 1510 -108
rect 1544 -142 1578 -108
rect 1612 -142 1646 -108
rect 1680 -142 1714 -108
rect 1748 -142 1856 -108
<< nsubdiff >>
rect 1402 1010 1498 1044
rect 1532 1010 1566 1044
rect 1600 1010 1634 1044
rect 1668 1010 1702 1044
rect 1736 1010 1770 1044
rect 1804 1010 1838 1044
rect 1872 1010 1906 1044
rect 1940 1010 1974 1044
rect 2008 1010 2042 1044
rect 2076 1010 2110 1044
rect 2144 1010 2240 1044
rect 1402 948 1436 1010
rect 2206 948 2240 1010
rect 1402 880 1436 914
rect 2206 880 2240 914
rect 1402 812 1436 846
rect 1402 744 1436 778
rect 1402 676 1436 710
rect 2206 812 2240 846
rect 2206 744 2240 778
rect 2206 676 2240 710
rect 1402 608 1436 642
rect 1402 512 1436 574
rect 2206 608 2240 642
rect 2206 512 2240 574
rect 1402 478 1498 512
rect 1532 478 1566 512
rect 1600 478 1634 512
rect 1668 478 1702 512
rect 1736 478 1770 512
rect 1804 478 1838 512
rect 1872 478 1906 512
rect 1940 478 1974 512
rect 2008 478 2042 512
rect 2076 478 2110 512
rect 2144 478 2240 512
<< psubdiffcont >>
rect 1510 372 1544 406
rect 1578 372 1612 406
rect 1646 372 1680 406
rect 1714 372 1748 406
rect 1402 251 1436 285
rect 1822 251 1856 285
rect 1402 183 1436 217
rect 1402 115 1436 149
rect 1402 47 1436 81
rect 1822 183 1856 217
rect 1822 115 1856 149
rect 1822 47 1856 81
rect 1402 -21 1436 13
rect 1822 -21 1856 13
rect 1510 -142 1544 -108
rect 1578 -142 1612 -108
rect 1646 -142 1680 -108
rect 1714 -142 1748 -108
<< nsubdiffcont >>
rect 1498 1010 1532 1044
rect 1566 1010 1600 1044
rect 1634 1010 1668 1044
rect 1702 1010 1736 1044
rect 1770 1010 1804 1044
rect 1838 1010 1872 1044
rect 1906 1010 1940 1044
rect 1974 1010 2008 1044
rect 2042 1010 2076 1044
rect 2110 1010 2144 1044
rect 1402 914 1436 948
rect 1402 846 1436 880
rect 2206 914 2240 948
rect 1402 778 1436 812
rect 1402 710 1436 744
rect 1402 642 1436 676
rect 2206 846 2240 880
rect 2206 778 2240 812
rect 2206 710 2240 744
rect 1402 574 1436 608
rect 2206 642 2240 676
rect 2206 574 2240 608
rect 1498 478 1532 512
rect 1566 478 1600 512
rect 1634 478 1668 512
rect 1702 478 1736 512
rect 1770 478 1804 512
rect 1838 478 1872 512
rect 1906 478 1940 512
rect 1974 478 2008 512
rect 2042 478 2076 512
rect 2110 478 2144 512
<< poly >>
rect 1566 886 2076 916
rect 1566 861 1596 886
rect 1662 861 1692 886
rect 1758 861 1788 886
rect 1854 861 1884 886
rect 1950 861 1980 886
rect 2046 861 2076 886
rect 1566 636 1596 661
rect 1662 636 1692 661
rect 1758 636 1788 661
rect 1854 636 1884 661
rect 1950 636 1980 661
rect 2046 636 2076 661
rect 1566 630 2076 636
rect 1548 614 2076 630
rect 1548 580 1564 614
rect 1598 606 1756 614
rect 1598 580 1614 606
rect 1548 564 1614 580
rect 1740 580 1756 606
rect 1790 606 1948 614
rect 1790 580 1806 606
rect 1740 564 1806 580
rect 1932 580 1948 606
rect 1982 606 2076 614
rect 1982 580 1998 606
rect 1932 564 1998 580
rect 1644 304 1710 320
rect 1644 284 1660 304
rect 1566 270 1660 284
rect 1694 270 1710 304
rect 1566 254 1710 270
rect 1566 232 1596 254
rect 1662 232 1692 254
rect 1566 10 1596 32
rect 1662 10 1692 32
rect 1566 -20 1692 10
<< polycont >>
rect 1564 580 1598 614
rect 1756 580 1790 614
rect 1948 580 1982 614
rect 1660 270 1694 304
<< locali >>
rect 1402 1010 1498 1044
rect 1532 1010 1566 1044
rect 1600 1010 1634 1044
rect 1668 1010 1702 1044
rect 1736 1010 1770 1044
rect 1402 948 1436 1010
rect 1402 880 1436 914
rect 1402 812 1436 846
rect 1402 744 1436 778
rect 1402 676 1436 710
rect 1516 846 1550 865
rect 1516 778 1550 780
rect 1516 742 1550 744
rect 1516 657 1550 676
rect 1612 846 1646 1010
rect 1612 778 1646 812
rect 1612 710 1646 744
rect 1612 657 1646 676
rect 1708 846 1742 865
rect 1708 778 1742 780
rect 1708 742 1742 744
rect 1708 657 1742 676
rect 1804 846 1838 1044
rect 1872 1010 1906 1044
rect 1940 1010 1974 1044
rect 2008 1010 2042 1044
rect 2076 1010 2110 1044
rect 2144 1010 2240 1044
rect 1804 778 1838 812
rect 1804 710 1838 744
rect 1804 657 1838 676
rect 1900 846 1934 865
rect 1900 778 1934 780
rect 1900 742 1934 744
rect 1900 657 1934 676
rect 1996 846 2030 1010
rect 2206 948 2240 1010
rect 2206 880 2240 914
rect 1996 778 2030 812
rect 1996 710 2030 744
rect 1996 657 2030 676
rect 2092 846 2126 865
rect 2092 778 2126 780
rect 2092 742 2126 744
rect 2092 657 2126 676
rect 2206 812 2240 846
rect 2206 744 2240 778
rect 2206 676 2240 710
rect 1402 608 1436 642
rect 1548 580 1564 614
rect 1598 580 1614 614
rect 1740 580 1756 614
rect 1790 580 1806 614
rect 1932 580 1948 614
rect 1982 580 1998 614
rect 2206 608 2240 642
rect 1402 512 1436 574
rect 2206 512 2240 574
rect 1402 478 1498 512
rect 1532 478 1566 512
rect 1600 478 1634 512
rect 1668 478 1702 512
rect 1736 478 1770 512
rect 1804 478 1838 512
rect 1872 478 1906 512
rect 1940 478 1974 512
rect 2008 478 2042 512
rect 2076 478 2110 512
rect 2144 478 2240 512
rect 1402 372 1510 406
rect 1544 372 1578 406
rect 1612 372 1646 406
rect 1680 372 1714 406
rect 1748 372 1856 406
rect 1402 285 1436 372
rect 1644 270 1660 304
rect 1694 270 1710 304
rect 1822 285 1856 372
rect 1402 217 1436 251
rect 1402 149 1436 183
rect 1402 81 1436 115
rect 1402 13 1436 47
rect 1516 217 1550 236
rect 1516 149 1550 151
rect 1516 113 1550 115
rect 1516 28 1550 47
rect 1612 217 1646 236
rect 1612 149 1646 183
rect 1612 81 1646 115
rect 1402 -108 1436 -21
rect 1402 -142 1510 -108
rect 1544 -142 1578 -108
rect 1612 -142 1646 47
rect 1708 217 1742 236
rect 1708 149 1742 151
rect 1708 113 1742 115
rect 1708 28 1742 47
rect 1822 217 1856 251
rect 1822 149 1856 183
rect 1822 81 1856 115
rect 1822 13 1856 47
rect 1822 -108 1856 -21
rect 1680 -142 1714 -108
rect 1748 -142 1856 -108
<< viali >>
rect 1516 812 1550 814
rect 1516 780 1550 812
rect 1516 710 1550 742
rect 1516 708 1550 710
rect 1708 812 1742 814
rect 1708 780 1742 812
rect 1708 710 1742 742
rect 1708 708 1742 710
rect 1900 812 1934 814
rect 1900 780 1934 812
rect 1900 710 1934 742
rect 1900 708 1934 710
rect 2092 812 2126 814
rect 2092 780 2126 812
rect 2092 710 2126 742
rect 2092 708 2126 710
rect 1564 580 1598 614
rect 1756 580 1790 614
rect 1948 580 1982 614
rect 1660 270 1694 304
rect 1516 183 1550 185
rect 1516 151 1550 183
rect 1516 81 1550 113
rect 1516 79 1550 81
rect 1708 183 1742 185
rect 1708 151 1742 183
rect 1708 81 1742 113
rect 1708 79 1742 81
<< metal1 >>
rect 1516 861 2126 876
rect 1510 848 2132 861
rect 1510 814 1556 848
rect 1510 780 1516 814
rect 1550 780 1556 814
rect 1510 742 1556 780
rect 1510 708 1516 742
rect 1550 708 1556 742
rect 1510 661 1556 708
rect 1702 814 1748 848
rect 1702 780 1708 814
rect 1742 780 1748 814
rect 1702 742 1748 780
rect 1702 708 1708 742
rect 1742 708 1748 742
rect 1702 661 1748 708
rect 1894 814 1940 848
rect 1894 780 1900 814
rect 1934 780 1940 814
rect 1894 742 1940 780
rect 1894 708 1900 742
rect 1934 708 1940 742
rect 1894 661 1940 708
rect 2086 814 2132 848
rect 2086 780 2092 814
rect 2126 780 2132 814
rect 2086 742 2132 780
rect 2086 708 2092 742
rect 2126 708 2132 742
rect 1552 614 1994 620
rect 1552 580 1564 614
rect 1598 580 1756 614
rect 1790 580 1948 614
rect 1982 580 1994 614
rect 1552 574 1994 580
rect 1660 310 1694 574
rect 2086 512 2132 708
rect 1822 478 2132 512
rect 1648 304 1706 310
rect 1648 270 1660 304
rect 1694 270 1706 304
rect 1648 264 1706 270
rect 1510 185 1556 232
rect 1510 151 1516 185
rect 1550 151 1556 185
rect 1510 113 1556 151
rect 1510 79 1516 113
rect 1550 79 1556 113
rect 1510 44 1556 79
rect 1702 185 1748 232
rect 1702 151 1708 185
rect 1742 151 1748 185
rect 1702 113 1748 151
rect 1702 79 1708 113
rect 1742 79 1748 113
rect 1702 44 1748 79
rect 1822 44 1856 478
rect 1510 32 1856 44
rect 1516 14 1856 32
<< labels >>
rlabel metal1 s 1674 432 1674 432 4 VIN
port 1 nsew
rlabel metal1 s 1838 430 1838 430 4 VOUT
port 2 nsew
rlabel locali s 2224 1024 2224 1024 4 VDD
port 3 nsew
rlabel locali s 1838 -122 1838 -122 4 VSS
port 4 nsew
<< end >>
