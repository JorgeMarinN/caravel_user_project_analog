magic
tech sky130A
magscale 1 2
timestamp 1640991954
<< locali >>
rect 5018 6437 5118 6470
rect 5018 6403 5051 6437
rect 5085 6403 5118 6437
rect 5018 6370 5118 6403
rect 4646 5225 4734 5252
rect 4646 5191 4673 5225
rect 4707 5191 4734 5225
rect 4646 5164 4734 5191
<< viali >>
rect 5051 6403 5085 6437
rect 4673 5191 4707 5225
<< metal1 >>
rect 5012 6437 5124 6476
rect 5012 6403 5051 6437
rect 5085 6403 5124 6437
rect 5012 6364 5124 6403
rect 3976 5666 4512 5784
rect 3976 5640 4144 5666
rect 3976 5524 4002 5640
rect 4118 5524 4144 5640
rect 3976 5498 4144 5524
rect 4674 5640 5310 5666
rect 4674 5524 5168 5640
rect 5284 5524 5310 5640
rect 4674 5498 5310 5524
rect 4634 5258 4744 5264
rect 6862 5258 6968 5264
rect 4634 5234 6968 5258
rect 4634 5225 6886 5234
rect 4634 5191 4673 5225
rect 4707 5191 6886 5225
rect 4634 5182 6886 5191
rect 6938 5182 6968 5234
rect 4634 5158 6968 5182
rect 4634 5152 4744 5158
rect 6862 5152 6968 5158
<< via1 >>
rect 4002 5524 4118 5640
rect 5168 5524 5284 5640
rect 6886 5182 6938 5234
<< metal2 >>
rect 3976 5640 4144 5666
rect 3976 5524 4002 5640
rect 4118 5524 4144 5640
rect 3976 5498 4144 5524
rect 5138 5650 5314 5670
rect 5138 5514 5158 5650
rect 5294 5514 5314 5650
rect 5138 5494 5314 5514
rect 6856 5234 6968 5264
rect 6856 5182 6886 5234
rect 6938 5182 6968 5234
rect 6856 5044 6968 5182
<< via2 >>
rect 5158 5640 5294 5650
rect 5158 5524 5168 5640
rect 5168 5524 5284 5640
rect 5284 5524 5294 5640
rect 5158 5514 5294 5524
<< metal3 >>
rect 5140 5654 5746 5666
rect 5140 5650 5590 5654
rect 5140 5514 5158 5650
rect 5294 5514 5590 5650
rect 5140 5510 5590 5514
rect 5734 5510 5746 5654
rect 5140 5498 5746 5510
<< via3 >>
rect 5590 5510 5734 5654
<< metal4 >>
rect 5584 5654 5740 5660
rect 5584 5510 5590 5654
rect 5734 5510 5740 5654
rect 5584 5504 5740 5510
use INV_v1p1  INV_v1p1_0
timestamp 1640991954
transform 1 0 2818 0 1 5366
box 1366 -168 2276 1080
use CAPOSC_v1p1  CAPOSC_v1p1_0
timestamp 1640991954
transform 1 0 -3068 0 1 432
box 3068 -432 10032 5306
<< labels >>
flabel metal3 s 5220 5580 5220 5580 0 FreeSans 2000 0 0 0 VOUT
port 1 nsew
flabel metal1 s 5034 6392 5034 6392 0 FreeSans 2000 0 0 0 VDD
port 2 nsew
flabel metal1 s 4984 5204 4984 5204 0 FreeSans 2000 0 0 0 VSS
port 3 nsew
<< end >>
